
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_Filter_Nb10_N11 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_Filter_Nb10_N11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Filter_Nb10_N11.all;

entity Filter_Nb10_N11 is

   port( DIN : in SIGNED (9 downto 0);  VIN, rst_n, clk : in std_logic;  B : in
         std_logic_vector (109 downto 0);  DOUT : out SIGNED (9 downto 0);  
         VOUT : out std_logic);

end Filter_Nb10_N11;

architecture SYN_beh of Filter_Nb10_N11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal x_vector_109_port, x_vector_108_port, x_vector_107_port, 
      x_vector_106_port, x_vector_105_port, x_vector_104_port, 
      x_vector_103_port, x_vector_102_port, x_vector_101_port, 
      x_vector_100_port, x_vector_99_port, x_vector_98_port, x_vector_97_port, 
      x_vector_96_port, x_vector_95_port, x_vector_94_port, x_vector_93_port, 
      x_vector_92_port, x_vector_91_port, x_vector_90_port, x_vector_89_port, 
      x_vector_88_port, x_vector_87_port, x_vector_86_port, x_vector_85_port, 
      x_vector_84_port, x_vector_83_port, x_vector_82_port, x_vector_81_port, 
      x_vector_80_port, x_vector_79_port, x_vector_78_port, x_vector_77_port, 
      x_vector_76_port, x_vector_75_port, x_vector_74_port, x_vector_73_port, 
      x_vector_72_port, x_vector_71_port, x_vector_70_port, x_vector_69_port, 
      x_vector_68_port, x_vector_67_port, x_vector_66_port, x_vector_65_port, 
      x_vector_64_port, x_vector_63_port, x_vector_62_port, x_vector_61_port, 
      x_vector_60_port, x_vector_59_port, x_vector_58_port, x_vector_57_port, 
      x_vector_56_port, x_vector_55_port, x_vector_54_port, x_vector_53_port, 
      x_vector_52_port, x_vector_51_port, x_vector_50_port, x_vector_49_port, 
      x_vector_48_port, x_vector_47_port, x_vector_46_port, x_vector_45_port, 
      x_vector_44_port, x_vector_43_port, x_vector_42_port, x_vector_41_port, 
      x_vector_40_port, x_vector_39_port, x_vector_38_port, x_vector_37_port, 
      x_vector_36_port, x_vector_35_port, x_vector_34_port, x_vector_33_port, 
      x_vector_32_port, x_vector_31_port, x_vector_30_port, x_vector_29_port, 
      x_vector_28_port, x_vector_27_port, x_vector_26_port, x_vector_25_port, 
      x_vector_24_port, x_vector_23_port, x_vector_22_port, x_vector_21_port, 
      x_vector_20_port, x_vector_19_port, x_vector_18_port, x_vector_17_port, 
      x_vector_16_port, x_vector_15_port, x_vector_14_port, x_vector_13_port, 
      x_vector_12_port, x_vector_11_port, x_vector_10_port, x_vector_9_port, 
      x_vector_8_port, x_vector_7_port, x_vector_6_port, x_vector_5_port, 
      x_vector_4_port, x_vector_3_port, x_vector_2_port, x_vector_1_port, 
      x_vector_0_port, N203, N204, N205, N206, N207, N208, N209, N210, N211, 
      N212, n21, n23, n72, n156, n157, n158, n159, n160, n161, n162, n163, n164
      , n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203_port, n204_port, n205_port, n206_port, n207_port, 
      n208_port, n209_port, n210_port, n211_port, n212_port, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N9, N89, N88, N87, N86,
      N85, N84, N83, N82, N81, N80, N8, N79, N78, N77, N76, N75, N74, N73, 
      N72_port, N71, N70, N7, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60,
      N6, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N5, N49, N48, N47, 
      N46, N45, N44, N43, N42, N41, N40, N4, N39, N38, N37, N36, N35, N34, N33,
      N32, N31, N30, N3, N29, N28, N27, N26, N25, N24, N23_port, N22, N21_port,
      N202_port, N201_port, N200_port, N20, N199_port, N198_port, N197_port, 
      N196_port, N195_port, N194_port, N193_port, N192_port, N191_port, 
      N190_port, N19, N189_port, N188_port, N187_port, N186_port, N185_port, 
      N184_port, N183_port, N182_port, N181_port, N180_port, N18, N179_port, 
      N178_port, N177_port, N176_port, N175_port, N174_port, N173_port, 
      N172_port, N171_port, N170_port, N17, N169_port, N168_port, N167_port, 
      N166_port, N165_port, N164_port, N163_port, N162_port, N161_port, 
      N160_port, N16, N159_port, N158_port, N157_port, N156_port, N155, N154, 
      N153, N152, N151, N150, N15, N149, N148, N147, N146, N145, N144, N143, 
      N142, N141, N140, N14, N139, N138, N137, N136, N135, N134, N133, N132, 
      N131, N130, N13, N129, N128, N127, N126, N125, N124, N123, N122, N121, 
      N120, N12, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
      N11, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N10, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, mult_42_n402, mult_42_n401, mult_42_n400, mult_42_n399, 
      mult_42_n398, mult_42_n397, mult_42_n396, mult_42_n395, mult_42_n394, 
      mult_42_n393, mult_42_n392, mult_42_n391, mult_42_n390, mult_42_n389, 
      mult_42_n388, mult_42_n387, mult_42_n386, mult_42_n385, mult_42_n384, 
      mult_42_n383, mult_42_n382, mult_42_n381, mult_42_n380, mult_42_n379, 
      mult_42_n378, mult_42_n377, mult_42_n376, mult_42_n375, mult_42_n374, 
      mult_42_n373, mult_42_n372, mult_42_n371, mult_42_n370, mult_42_n369, 
      mult_42_n368, mult_42_n367, mult_42_n366, mult_42_n365, mult_42_n364, 
      mult_42_n363, mult_42_n362, mult_42_n361, mult_42_n360, mult_42_n359, 
      mult_42_n358, mult_42_n357, mult_42_n356, mult_42_n355, mult_42_n354, 
      mult_42_n353, mult_42_n352, mult_42_n351, mult_42_n350, mult_42_n349, 
      mult_42_n348, mult_42_n347, mult_42_n346, mult_42_n345, mult_42_n344, 
      mult_42_n343, mult_42_n342, mult_42_n341, mult_42_n340, mult_42_n339, 
      mult_42_n338, mult_42_n337, mult_42_n336, mult_42_n335, mult_42_n334, 
      mult_42_n333, mult_42_n332, mult_42_n331, mult_42_n330, mult_42_n329, 
      mult_42_n328, mult_42_n327, mult_42_n326, mult_42_n325, mult_42_n324, 
      mult_42_n323, mult_42_n322, mult_42_n321, mult_42_n320, mult_42_n319, 
      mult_42_n318, mult_42_n317, mult_42_n316, mult_42_n315, mult_42_n314, 
      mult_42_n313, mult_42_n312, mult_42_n311, mult_42_n310, mult_42_n309, 
      mult_42_n308, mult_42_n307, mult_42_n306, mult_42_n305, mult_42_n304, 
      mult_42_n303, mult_42_n302, mult_42_n301, mult_42_n300, mult_42_n299, 
      mult_42_n298, mult_42_n297, mult_42_n296, mult_42_n295, mult_42_n157, 
      mult_42_n156, mult_42_n155, mult_42_n154, mult_42_n153, mult_42_n152, 
      mult_42_n151, mult_42_n148, mult_42_n147, mult_42_n146, mult_42_n145, 
      mult_42_n144, mult_42_n143, mult_42_n142, mult_42_n140, mult_42_n139, 
      mult_42_n138, mult_42_n137, mult_42_n136, mult_42_n135, mult_42_n134, 
      mult_42_n133, mult_42_n132, mult_42_n131, mult_42_n129, mult_42_n128, 
      mult_42_n127, mult_42_n126, mult_42_n124, mult_42_n123, mult_42_n122, 
      mult_42_n121, mult_42_n119, mult_42_n118, mult_42_n117, mult_42_n116, 
      mult_42_n115, mult_42_n114, mult_42_n113, mult_42_n112, mult_42_n111, 
      mult_42_n107, mult_42_n106, mult_42_n105, mult_42_n90, mult_42_n89, 
      mult_42_n88, mult_42_n87, mult_42_n86, mult_42_n85, mult_42_n84, 
      mult_42_n83, mult_42_n82, mult_42_n81, mult_42_n80, mult_42_n79, 
      mult_42_n78, mult_42_n77, mult_42_n76, mult_42_n75, mult_42_n74, 
      mult_42_n73, mult_42_n72, mult_42_n71, mult_42_n70, mult_42_n69, 
      mult_42_n68, mult_42_n67, mult_42_n66, mult_42_n65, mult_42_n64, 
      mult_42_n63, mult_42_n62, mult_42_n61, mult_42_n60, mult_42_n59, 
      mult_42_n58, mult_42_n57, mult_42_n56, mult_42_n55, mult_42_n54, 
      mult_42_n53, mult_42_n52, mult_42_n51, mult_42_n50, mult_42_n48, 
      mult_42_n47, mult_42_n46, mult_42_n45, mult_42_n44, mult_42_n43, 
      mult_42_n42, mult_42_n41, mult_42_n40, mult_42_n39, mult_42_n38, 
      mult_42_n37, mult_42_n35, mult_42_n34, mult_42_n33, mult_42_n32, 
      mult_42_n31, mult_42_n30, mult_42_n29, mult_42_n28, mult_42_n27, 
      mult_42_n25, mult_42_n24, mult_42_n23, mult_42_n22, mult_42_n21, 
      mult_42_n19, mult_42_n10, mult_42_n9, mult_42_n8, mult_42_n7, mult_42_n6,
      mult_42_n5, mult_42_n4, mult_42_n3, mult_42_n2, mult_42_n1, 
      mult_42_I2_n402, mult_42_I2_n401, mult_42_I2_n400, mult_42_I2_n399, 
      mult_42_I2_n398, mult_42_I2_n397, mult_42_I2_n396, mult_42_I2_n395, 
      mult_42_I2_n394, mult_42_I2_n393, mult_42_I2_n392, mult_42_I2_n391, 
      mult_42_I2_n390, mult_42_I2_n389, mult_42_I2_n388, mult_42_I2_n387, 
      mult_42_I2_n386, mult_42_I2_n385, mult_42_I2_n384, mult_42_I2_n383, 
      mult_42_I2_n382, mult_42_I2_n381, mult_42_I2_n380, mult_42_I2_n379, 
      mult_42_I2_n378, mult_42_I2_n377, mult_42_I2_n376, mult_42_I2_n375, 
      mult_42_I2_n374, mult_42_I2_n373, mult_42_I2_n372, mult_42_I2_n371, 
      mult_42_I2_n370, mult_42_I2_n369, mult_42_I2_n368, mult_42_I2_n367, 
      mult_42_I2_n366, mult_42_I2_n365, mult_42_I2_n364, mult_42_I2_n363, 
      mult_42_I2_n362, mult_42_I2_n361, mult_42_I2_n360, mult_42_I2_n359, 
      mult_42_I2_n358, mult_42_I2_n357, mult_42_I2_n356, mult_42_I2_n355, 
      mult_42_I2_n354, mult_42_I2_n353, mult_42_I2_n352, mult_42_I2_n351, 
      mult_42_I2_n350, mult_42_I2_n349, mult_42_I2_n348, mult_42_I2_n347, 
      mult_42_I2_n346, mult_42_I2_n345, mult_42_I2_n344, mult_42_I2_n343, 
      mult_42_I2_n342, mult_42_I2_n341, mult_42_I2_n340, mult_42_I2_n339, 
      mult_42_I2_n338, mult_42_I2_n337, mult_42_I2_n336, mult_42_I2_n335, 
      mult_42_I2_n334, mult_42_I2_n333, mult_42_I2_n332, mult_42_I2_n331, 
      mult_42_I2_n330, mult_42_I2_n329, mult_42_I2_n328, mult_42_I2_n327, 
      mult_42_I2_n326, mult_42_I2_n325, mult_42_I2_n324, mult_42_I2_n323, 
      mult_42_I2_n322, mult_42_I2_n321, mult_42_I2_n320, mult_42_I2_n319, 
      mult_42_I2_n318, mult_42_I2_n317, mult_42_I2_n316, mult_42_I2_n315, 
      mult_42_I2_n314, mult_42_I2_n313, mult_42_I2_n312, mult_42_I2_n311, 
      mult_42_I2_n310, mult_42_I2_n309, mult_42_I2_n308, mult_42_I2_n307, 
      mult_42_I2_n306, mult_42_I2_n305, mult_42_I2_n304, mult_42_I2_n303, 
      mult_42_I2_n302, mult_42_I2_n301, mult_42_I2_n300, mult_42_I2_n299, 
      mult_42_I2_n298, mult_42_I2_n297, mult_42_I2_n296, mult_42_I2_n295, 
      mult_42_I2_n157, mult_42_I2_n156, mult_42_I2_n155, mult_42_I2_n154, 
      mult_42_I2_n153, mult_42_I2_n152, mult_42_I2_n151, mult_42_I2_n148, 
      mult_42_I2_n147, mult_42_I2_n146, mult_42_I2_n145, mult_42_I2_n144, 
      mult_42_I2_n143, mult_42_I2_n142, mult_42_I2_n140, mult_42_I2_n139, 
      mult_42_I2_n138, mult_42_I2_n137, mult_42_I2_n136, mult_42_I2_n135, 
      mult_42_I2_n134, mult_42_I2_n133, mult_42_I2_n132, mult_42_I2_n131, 
      mult_42_I2_n129, mult_42_I2_n128, mult_42_I2_n127, mult_42_I2_n126, 
      mult_42_I2_n124, mult_42_I2_n123, mult_42_I2_n122, mult_42_I2_n121, 
      mult_42_I2_n119, mult_42_I2_n118, mult_42_I2_n117, mult_42_I2_n116, 
      mult_42_I2_n115, mult_42_I2_n114, mult_42_I2_n113, mult_42_I2_n112, 
      mult_42_I2_n111, mult_42_I2_n107, mult_42_I2_n106, mult_42_I2_n105, 
      mult_42_I2_n90, mult_42_I2_n89, mult_42_I2_n88, mult_42_I2_n87, 
      mult_42_I2_n86, mult_42_I2_n85, mult_42_I2_n84, mult_42_I2_n83, 
      mult_42_I2_n82, mult_42_I2_n81, mult_42_I2_n80, mult_42_I2_n79, 
      mult_42_I2_n78, mult_42_I2_n77, mult_42_I2_n76, mult_42_I2_n75, 
      mult_42_I2_n74, mult_42_I2_n73, mult_42_I2_n72, mult_42_I2_n71, 
      mult_42_I2_n70, mult_42_I2_n69, mult_42_I2_n68, mult_42_I2_n67, 
      mult_42_I2_n66, mult_42_I2_n65, mult_42_I2_n64, mult_42_I2_n63, 
      mult_42_I2_n62, mult_42_I2_n61, mult_42_I2_n60, mult_42_I2_n59, 
      mult_42_I2_n58, mult_42_I2_n57, mult_42_I2_n56, mult_42_I2_n55, 
      mult_42_I2_n54, mult_42_I2_n53, mult_42_I2_n52, mult_42_I2_n51, 
      mult_42_I2_n50, mult_42_I2_n48, mult_42_I2_n47, mult_42_I2_n46, 
      mult_42_I2_n45, mult_42_I2_n44, mult_42_I2_n43, mult_42_I2_n42, 
      mult_42_I2_n41, mult_42_I2_n40, mult_42_I2_n39, mult_42_I2_n38, 
      mult_42_I2_n37, mult_42_I2_n35, mult_42_I2_n34, mult_42_I2_n33, 
      mult_42_I2_n32, mult_42_I2_n31, mult_42_I2_n30, mult_42_I2_n29, 
      mult_42_I2_n28, mult_42_I2_n27, mult_42_I2_n25, mult_42_I2_n24, 
      mult_42_I2_n23, mult_42_I2_n22, mult_42_I2_n21, mult_42_I2_n19, 
      mult_42_I2_n10, mult_42_I2_n9, mult_42_I2_n8, mult_42_I2_n7, 
      mult_42_I2_n6, mult_42_I2_n5, mult_42_I2_n4, mult_42_I2_n3, mult_42_I2_n2
      , mult_42_I2_n1, mult_42_I3_n402, mult_42_I3_n401, mult_42_I3_n400, 
      mult_42_I3_n399, mult_42_I3_n398, mult_42_I3_n397, mult_42_I3_n396, 
      mult_42_I3_n395, mult_42_I3_n394, mult_42_I3_n393, mult_42_I3_n392, 
      mult_42_I3_n391, mult_42_I3_n390, mult_42_I3_n389, mult_42_I3_n388, 
      mult_42_I3_n387, mult_42_I3_n386, mult_42_I3_n385, mult_42_I3_n384, 
      mult_42_I3_n383, mult_42_I3_n382, mult_42_I3_n381, mult_42_I3_n380, 
      mult_42_I3_n379, mult_42_I3_n378, mult_42_I3_n377, mult_42_I3_n376, 
      mult_42_I3_n375, mult_42_I3_n374, mult_42_I3_n373, mult_42_I3_n372, 
      mult_42_I3_n371, mult_42_I3_n370, mult_42_I3_n369, mult_42_I3_n368, 
      mult_42_I3_n367, mult_42_I3_n366, mult_42_I3_n365, mult_42_I3_n364, 
      mult_42_I3_n363, mult_42_I3_n362, mult_42_I3_n361, mult_42_I3_n360, 
      mult_42_I3_n359, mult_42_I3_n358, mult_42_I3_n357, mult_42_I3_n356, 
      mult_42_I3_n355, mult_42_I3_n354, mult_42_I3_n353, mult_42_I3_n352, 
      mult_42_I3_n351, mult_42_I3_n350, mult_42_I3_n349, mult_42_I3_n348, 
      mult_42_I3_n347, mult_42_I3_n346, mult_42_I3_n345, mult_42_I3_n344, 
      mult_42_I3_n343, mult_42_I3_n342, mult_42_I3_n341, mult_42_I3_n340, 
      mult_42_I3_n339, mult_42_I3_n338, mult_42_I3_n337, mult_42_I3_n336, 
      mult_42_I3_n335, mult_42_I3_n334, mult_42_I3_n333, mult_42_I3_n332, 
      mult_42_I3_n331, mult_42_I3_n330, mult_42_I3_n329, mult_42_I3_n328, 
      mult_42_I3_n327, mult_42_I3_n326, mult_42_I3_n325, mult_42_I3_n324, 
      mult_42_I3_n323, mult_42_I3_n322, mult_42_I3_n321, mult_42_I3_n320, 
      mult_42_I3_n319, mult_42_I3_n318, mult_42_I3_n317, mult_42_I3_n316, 
      mult_42_I3_n315, mult_42_I3_n314, mult_42_I3_n313, mult_42_I3_n312, 
      mult_42_I3_n311, mult_42_I3_n310, mult_42_I3_n309, mult_42_I3_n308, 
      mult_42_I3_n307, mult_42_I3_n306, mult_42_I3_n305, mult_42_I3_n304, 
      mult_42_I3_n303, mult_42_I3_n302, mult_42_I3_n301, mult_42_I3_n300, 
      mult_42_I3_n299, mult_42_I3_n298, mult_42_I3_n297, mult_42_I3_n296, 
      mult_42_I3_n295, mult_42_I3_n157, mult_42_I3_n156, mult_42_I3_n155, 
      mult_42_I3_n154, mult_42_I3_n153, mult_42_I3_n152, mult_42_I3_n151, 
      mult_42_I3_n148, mult_42_I3_n147, mult_42_I3_n146, mult_42_I3_n145, 
      mult_42_I3_n144, mult_42_I3_n143, mult_42_I3_n142, mult_42_I3_n140, 
      mult_42_I3_n139, mult_42_I3_n138, mult_42_I3_n137, mult_42_I3_n136, 
      mult_42_I3_n135, mult_42_I3_n134, mult_42_I3_n133, mult_42_I3_n132, 
      mult_42_I3_n131, mult_42_I3_n129, mult_42_I3_n128, mult_42_I3_n127, 
      mult_42_I3_n126, mult_42_I3_n124, mult_42_I3_n123, mult_42_I3_n122, 
      mult_42_I3_n121, mult_42_I3_n119, mult_42_I3_n118, mult_42_I3_n117, 
      mult_42_I3_n116, mult_42_I3_n115, mult_42_I3_n114, mult_42_I3_n113, 
      mult_42_I3_n112, mult_42_I3_n111, mult_42_I3_n107, mult_42_I3_n106, 
      mult_42_I3_n105, mult_42_I3_n90, mult_42_I3_n89, mult_42_I3_n88, 
      mult_42_I3_n87, mult_42_I3_n86, mult_42_I3_n85, mult_42_I3_n84, 
      mult_42_I3_n83, mult_42_I3_n82, mult_42_I3_n81, mult_42_I3_n80, 
      mult_42_I3_n79, mult_42_I3_n78, mult_42_I3_n77, mult_42_I3_n76, 
      mult_42_I3_n75, mult_42_I3_n74, mult_42_I3_n73, mult_42_I3_n72, 
      mult_42_I3_n71, mult_42_I3_n70, mult_42_I3_n69, mult_42_I3_n68, 
      mult_42_I3_n67, mult_42_I3_n66, mult_42_I3_n65, mult_42_I3_n64, 
      mult_42_I3_n63, mult_42_I3_n62, mult_42_I3_n61, mult_42_I3_n60, 
      mult_42_I3_n59, mult_42_I3_n58, mult_42_I3_n57, mult_42_I3_n56, 
      mult_42_I3_n55, mult_42_I3_n54, mult_42_I3_n53, mult_42_I3_n52, 
      mult_42_I3_n51, mult_42_I3_n50, mult_42_I3_n48, mult_42_I3_n47, 
      mult_42_I3_n46, mult_42_I3_n45, mult_42_I3_n44, mult_42_I3_n43, 
      mult_42_I3_n42, mult_42_I3_n41, mult_42_I3_n40, mult_42_I3_n39, 
      mult_42_I3_n38, mult_42_I3_n37, mult_42_I3_n35, mult_42_I3_n34, 
      mult_42_I3_n33, mult_42_I3_n32, mult_42_I3_n31, mult_42_I3_n30, 
      mult_42_I3_n29, mult_42_I3_n28, mult_42_I3_n27, mult_42_I3_n25, 
      mult_42_I3_n24, mult_42_I3_n23, mult_42_I3_n22, mult_42_I3_n21, 
      mult_42_I3_n19, mult_42_I3_n10, mult_42_I3_n9, mult_42_I3_n8, 
      mult_42_I3_n7, mult_42_I3_n6, mult_42_I3_n5, mult_42_I3_n4, mult_42_I3_n3
      , mult_42_I3_n2, mult_42_I3_n1, mult_42_I4_n402, mult_42_I4_n401, 
      mult_42_I4_n400, mult_42_I4_n399, mult_42_I4_n398, mult_42_I4_n397, 
      mult_42_I4_n396, mult_42_I4_n395, mult_42_I4_n394, mult_42_I4_n393, 
      mult_42_I4_n392, mult_42_I4_n391, mult_42_I4_n390, mult_42_I4_n389, 
      mult_42_I4_n388, mult_42_I4_n387, mult_42_I4_n386, mult_42_I4_n385, 
      mult_42_I4_n384, mult_42_I4_n383, mult_42_I4_n382, mult_42_I4_n381, 
      mult_42_I4_n380, mult_42_I4_n379, mult_42_I4_n378, mult_42_I4_n377, 
      mult_42_I4_n376, mult_42_I4_n375, mult_42_I4_n374, mult_42_I4_n373, 
      mult_42_I4_n372, mult_42_I4_n371, mult_42_I4_n370, mult_42_I4_n369, 
      mult_42_I4_n368, mult_42_I4_n367, mult_42_I4_n366, mult_42_I4_n365, 
      mult_42_I4_n364, mult_42_I4_n363, mult_42_I4_n362, mult_42_I4_n361, 
      mult_42_I4_n360, mult_42_I4_n359, mult_42_I4_n358, mult_42_I4_n357, 
      mult_42_I4_n356, mult_42_I4_n355, mult_42_I4_n354, mult_42_I4_n353, 
      mult_42_I4_n352, mult_42_I4_n351, mult_42_I4_n350, mult_42_I4_n349, 
      mult_42_I4_n348, mult_42_I4_n347, mult_42_I4_n346, mult_42_I4_n345, 
      mult_42_I4_n344, mult_42_I4_n343, mult_42_I4_n342, mult_42_I4_n341, 
      mult_42_I4_n340, mult_42_I4_n339, mult_42_I4_n338, mult_42_I4_n337, 
      mult_42_I4_n336, mult_42_I4_n335, mult_42_I4_n334, mult_42_I4_n333, 
      mult_42_I4_n332, mult_42_I4_n331, mult_42_I4_n330, mult_42_I4_n329, 
      mult_42_I4_n328, mult_42_I4_n327, mult_42_I4_n326, mult_42_I4_n325, 
      mult_42_I4_n324, mult_42_I4_n323, mult_42_I4_n322, mult_42_I4_n321, 
      mult_42_I4_n320, mult_42_I4_n319, mult_42_I4_n318, mult_42_I4_n317, 
      mult_42_I4_n316, mult_42_I4_n315, mult_42_I4_n314, mult_42_I4_n313, 
      mult_42_I4_n312, mult_42_I4_n311, mult_42_I4_n310, mult_42_I4_n309, 
      mult_42_I4_n308, mult_42_I4_n307, mult_42_I4_n306, mult_42_I4_n305, 
      mult_42_I4_n304, mult_42_I4_n303, mult_42_I4_n302, mult_42_I4_n301, 
      mult_42_I4_n300, mult_42_I4_n299, mult_42_I4_n298, mult_42_I4_n297, 
      mult_42_I4_n296, mult_42_I4_n295, mult_42_I4_n157, mult_42_I4_n156, 
      mult_42_I4_n155, mult_42_I4_n154, mult_42_I4_n153, mult_42_I4_n152, 
      mult_42_I4_n151, mult_42_I4_n148, mult_42_I4_n147, mult_42_I4_n146, 
      mult_42_I4_n145, mult_42_I4_n144, mult_42_I4_n143, mult_42_I4_n142, 
      mult_42_I4_n140, mult_42_I4_n139, mult_42_I4_n138, mult_42_I4_n137, 
      mult_42_I4_n136, mult_42_I4_n135, mult_42_I4_n134, mult_42_I4_n133, 
      mult_42_I4_n132, mult_42_I4_n131, mult_42_I4_n129, mult_42_I4_n128, 
      mult_42_I4_n127, mult_42_I4_n126, mult_42_I4_n124, mult_42_I4_n123, 
      mult_42_I4_n122, mult_42_I4_n121, mult_42_I4_n119, mult_42_I4_n118, 
      mult_42_I4_n117, mult_42_I4_n116, mult_42_I4_n115, mult_42_I4_n114, 
      mult_42_I4_n113, mult_42_I4_n112, mult_42_I4_n111, mult_42_I4_n107, 
      mult_42_I4_n106, mult_42_I4_n105, mult_42_I4_n90, mult_42_I4_n89, 
      mult_42_I4_n88, mult_42_I4_n87, mult_42_I4_n86, mult_42_I4_n85, 
      mult_42_I4_n84, mult_42_I4_n83, mult_42_I4_n82, mult_42_I4_n81, 
      mult_42_I4_n80, mult_42_I4_n79, mult_42_I4_n78, mult_42_I4_n77, 
      mult_42_I4_n76, mult_42_I4_n75, mult_42_I4_n74, mult_42_I4_n73, 
      mult_42_I4_n72, mult_42_I4_n71, mult_42_I4_n70, mult_42_I4_n69, 
      mult_42_I4_n68, mult_42_I4_n67, mult_42_I4_n66, mult_42_I4_n65, 
      mult_42_I4_n64, mult_42_I4_n63, mult_42_I4_n62, mult_42_I4_n61, 
      mult_42_I4_n60, mult_42_I4_n59, mult_42_I4_n58, mult_42_I4_n57, 
      mult_42_I4_n56, mult_42_I4_n55, mult_42_I4_n54, mult_42_I4_n53, 
      mult_42_I4_n52, mult_42_I4_n51, mult_42_I4_n50, mult_42_I4_n48, 
      mult_42_I4_n47, mult_42_I4_n46, mult_42_I4_n45, mult_42_I4_n44, 
      mult_42_I4_n43, mult_42_I4_n42, mult_42_I4_n41, mult_42_I4_n40, 
      mult_42_I4_n39, mult_42_I4_n38, mult_42_I4_n37, mult_42_I4_n35, 
      mult_42_I4_n34, mult_42_I4_n33, mult_42_I4_n32, mult_42_I4_n31, 
      mult_42_I4_n30, mult_42_I4_n29, mult_42_I4_n28, mult_42_I4_n27, 
      mult_42_I4_n25, mult_42_I4_n24, mult_42_I4_n23, mult_42_I4_n22, 
      mult_42_I4_n21, mult_42_I4_n19, mult_42_I4_n10, mult_42_I4_n9, 
      mult_42_I4_n8, mult_42_I4_n7, mult_42_I4_n6, mult_42_I4_n5, mult_42_I4_n4
      , mult_42_I4_n3, mult_42_I4_n2, mult_42_I4_n1, mult_42_I5_n402, 
      mult_42_I5_n401, mult_42_I5_n400, mult_42_I5_n399, mult_42_I5_n398, 
      mult_42_I5_n397, mult_42_I5_n396, mult_42_I5_n395, mult_42_I5_n394, 
      mult_42_I5_n393, mult_42_I5_n392, mult_42_I5_n391, mult_42_I5_n390, 
      mult_42_I5_n389, mult_42_I5_n388, mult_42_I5_n387, mult_42_I5_n386, 
      mult_42_I5_n385, mult_42_I5_n384, mult_42_I5_n383, mult_42_I5_n382, 
      mult_42_I5_n381, mult_42_I5_n380, mult_42_I5_n379, mult_42_I5_n378, 
      mult_42_I5_n377, mult_42_I5_n376, mult_42_I5_n375, mult_42_I5_n374, 
      mult_42_I5_n373, mult_42_I5_n372, mult_42_I5_n371, mult_42_I5_n370, 
      mult_42_I5_n369, mult_42_I5_n368, mult_42_I5_n367, mult_42_I5_n366, 
      mult_42_I5_n365, mult_42_I5_n364, mult_42_I5_n363, mult_42_I5_n362, 
      mult_42_I5_n361, mult_42_I5_n360, mult_42_I5_n359, mult_42_I5_n358, 
      mult_42_I5_n357, mult_42_I5_n356, mult_42_I5_n355, mult_42_I5_n354, 
      mult_42_I5_n353, mult_42_I5_n352, mult_42_I5_n351, mult_42_I5_n350, 
      mult_42_I5_n349, mult_42_I5_n348, mult_42_I5_n347, mult_42_I5_n346, 
      mult_42_I5_n345, mult_42_I5_n344, mult_42_I5_n343, mult_42_I5_n342, 
      mult_42_I5_n341, mult_42_I5_n340, mult_42_I5_n339, mult_42_I5_n338, 
      mult_42_I5_n337, mult_42_I5_n336, mult_42_I5_n335, mult_42_I5_n334, 
      mult_42_I5_n333, mult_42_I5_n332, mult_42_I5_n331, mult_42_I5_n330, 
      mult_42_I5_n329, mult_42_I5_n328, mult_42_I5_n327, mult_42_I5_n326, 
      mult_42_I5_n325, mult_42_I5_n324, mult_42_I5_n323, mult_42_I5_n322, 
      mult_42_I5_n321, mult_42_I5_n320, mult_42_I5_n319, mult_42_I5_n318, 
      mult_42_I5_n317, mult_42_I5_n316, mult_42_I5_n315, mult_42_I5_n314, 
      mult_42_I5_n313, mult_42_I5_n312, mult_42_I5_n311, mult_42_I5_n310, 
      mult_42_I5_n309, mult_42_I5_n308, mult_42_I5_n307, mult_42_I5_n306, 
      mult_42_I5_n305, mult_42_I5_n304, mult_42_I5_n303, mult_42_I5_n302, 
      mult_42_I5_n301, mult_42_I5_n300, mult_42_I5_n299, mult_42_I5_n298, 
      mult_42_I5_n297, mult_42_I5_n296, mult_42_I5_n295, mult_42_I5_n157, 
      mult_42_I5_n156, mult_42_I5_n155, mult_42_I5_n154, mult_42_I5_n153, 
      mult_42_I5_n152, mult_42_I5_n151, mult_42_I5_n148, mult_42_I5_n147, 
      mult_42_I5_n146, mult_42_I5_n145, mult_42_I5_n144, mult_42_I5_n143, 
      mult_42_I5_n142, mult_42_I5_n140, mult_42_I5_n139, mult_42_I5_n138, 
      mult_42_I5_n137, mult_42_I5_n136, mult_42_I5_n135, mult_42_I5_n134, 
      mult_42_I5_n133, mult_42_I5_n132, mult_42_I5_n131, mult_42_I5_n129, 
      mult_42_I5_n128, mult_42_I5_n127, mult_42_I5_n126, mult_42_I5_n124, 
      mult_42_I5_n123, mult_42_I5_n122, mult_42_I5_n121, mult_42_I5_n119, 
      mult_42_I5_n118, mult_42_I5_n117, mult_42_I5_n116, mult_42_I5_n115, 
      mult_42_I5_n114, mult_42_I5_n113, mult_42_I5_n112, mult_42_I5_n111, 
      mult_42_I5_n107, mult_42_I5_n106, mult_42_I5_n105, mult_42_I5_n90, 
      mult_42_I5_n89, mult_42_I5_n88, mult_42_I5_n87, mult_42_I5_n86, 
      mult_42_I5_n85, mult_42_I5_n84, mult_42_I5_n83, mult_42_I5_n82, 
      mult_42_I5_n81, mult_42_I5_n80, mult_42_I5_n79, mult_42_I5_n78, 
      mult_42_I5_n77, mult_42_I5_n76, mult_42_I5_n75, mult_42_I5_n74, 
      mult_42_I5_n73, mult_42_I5_n72, mult_42_I5_n71, mult_42_I5_n70, 
      mult_42_I5_n69, mult_42_I5_n68, mult_42_I5_n67, mult_42_I5_n66, 
      mult_42_I5_n65, mult_42_I5_n64, mult_42_I5_n63, mult_42_I5_n62, 
      mult_42_I5_n61, mult_42_I5_n60, mult_42_I5_n59, mult_42_I5_n58, 
      mult_42_I5_n57, mult_42_I5_n56, mult_42_I5_n55, mult_42_I5_n54, 
      mult_42_I5_n53, mult_42_I5_n52, mult_42_I5_n51, mult_42_I5_n50, 
      mult_42_I5_n48, mult_42_I5_n47, mult_42_I5_n46, mult_42_I5_n45, 
      mult_42_I5_n44, mult_42_I5_n43, mult_42_I5_n42, mult_42_I5_n41, 
      mult_42_I5_n40, mult_42_I5_n39, mult_42_I5_n38, mult_42_I5_n37, 
      mult_42_I5_n35, mult_42_I5_n34, mult_42_I5_n33, mult_42_I5_n32, 
      mult_42_I5_n31, mult_42_I5_n30, mult_42_I5_n29, mult_42_I5_n28, 
      mult_42_I5_n27, mult_42_I5_n25, mult_42_I5_n24, mult_42_I5_n23, 
      mult_42_I5_n22, mult_42_I5_n21, mult_42_I5_n19, mult_42_I5_n10, 
      mult_42_I5_n9, mult_42_I5_n8, mult_42_I5_n7, mult_42_I5_n6, mult_42_I5_n5
      , mult_42_I5_n4, mult_42_I5_n3, mult_42_I5_n2, mult_42_I5_n1, 
      mult_42_I6_n402, mult_42_I6_n401, mult_42_I6_n400, mult_42_I6_n399, 
      mult_42_I6_n398, mult_42_I6_n397, mult_42_I6_n396, mult_42_I6_n395, 
      mult_42_I6_n394, mult_42_I6_n393, mult_42_I6_n392, mult_42_I6_n391, 
      mult_42_I6_n390, mult_42_I6_n389, mult_42_I6_n388, mult_42_I6_n387, 
      mult_42_I6_n386, mult_42_I6_n385, mult_42_I6_n384, mult_42_I6_n383, 
      mult_42_I6_n382, mult_42_I6_n381, mult_42_I6_n380, mult_42_I6_n379, 
      mult_42_I6_n378, mult_42_I6_n377, mult_42_I6_n376, mult_42_I6_n375, 
      mult_42_I6_n374, mult_42_I6_n373, mult_42_I6_n372, mult_42_I6_n371, 
      mult_42_I6_n370, mult_42_I6_n369, mult_42_I6_n368, mult_42_I6_n367, 
      mult_42_I6_n366, mult_42_I6_n365, mult_42_I6_n364, mult_42_I6_n363, 
      mult_42_I6_n362, mult_42_I6_n361, mult_42_I6_n360, mult_42_I6_n359, 
      mult_42_I6_n358, mult_42_I6_n357, mult_42_I6_n356, mult_42_I6_n355, 
      mult_42_I6_n354, mult_42_I6_n353, mult_42_I6_n352, mult_42_I6_n351, 
      mult_42_I6_n350, mult_42_I6_n349, mult_42_I6_n348, mult_42_I6_n347, 
      mult_42_I6_n346, mult_42_I6_n345, mult_42_I6_n344, mult_42_I6_n343, 
      mult_42_I6_n342, mult_42_I6_n341, mult_42_I6_n340, mult_42_I6_n339, 
      mult_42_I6_n338, mult_42_I6_n337, mult_42_I6_n336, mult_42_I6_n335, 
      mult_42_I6_n334, mult_42_I6_n333, mult_42_I6_n332, mult_42_I6_n331, 
      mult_42_I6_n330, mult_42_I6_n329, mult_42_I6_n328, mult_42_I6_n327, 
      mult_42_I6_n326, mult_42_I6_n325, mult_42_I6_n324, mult_42_I6_n323, 
      mult_42_I6_n322, mult_42_I6_n321, mult_42_I6_n320, mult_42_I6_n319, 
      mult_42_I6_n318, mult_42_I6_n317, mult_42_I6_n316, mult_42_I6_n315, 
      mult_42_I6_n314, mult_42_I6_n313, mult_42_I6_n312, mult_42_I6_n311, 
      mult_42_I6_n310, mult_42_I6_n309, mult_42_I6_n308, mult_42_I6_n307, 
      mult_42_I6_n306, mult_42_I6_n305, mult_42_I6_n304, mult_42_I6_n303, 
      mult_42_I6_n302, mult_42_I6_n301, mult_42_I6_n300, mult_42_I6_n299, 
      mult_42_I6_n298, mult_42_I6_n297, mult_42_I6_n296, mult_42_I6_n295, 
      mult_42_I6_n157, mult_42_I6_n156, mult_42_I6_n155, mult_42_I6_n154, 
      mult_42_I6_n153, mult_42_I6_n152, mult_42_I6_n151, mult_42_I6_n148, 
      mult_42_I6_n147, mult_42_I6_n146, mult_42_I6_n145, mult_42_I6_n144, 
      mult_42_I6_n143, mult_42_I6_n142, mult_42_I6_n140, mult_42_I6_n139, 
      mult_42_I6_n138, mult_42_I6_n137, mult_42_I6_n136, mult_42_I6_n135, 
      mult_42_I6_n134, mult_42_I6_n133, mult_42_I6_n132, mult_42_I6_n131, 
      mult_42_I6_n129, mult_42_I6_n128, mult_42_I6_n127, mult_42_I6_n126, 
      mult_42_I6_n124, mult_42_I6_n123, mult_42_I6_n122, mult_42_I6_n121, 
      mult_42_I6_n119, mult_42_I6_n118, mult_42_I6_n117, mult_42_I6_n116, 
      mult_42_I6_n115, mult_42_I6_n114, mult_42_I6_n113, mult_42_I6_n112, 
      mult_42_I6_n111, mult_42_I6_n107, mult_42_I6_n106, mult_42_I6_n105, 
      mult_42_I6_n90, mult_42_I6_n89, mult_42_I6_n88, mult_42_I6_n87, 
      mult_42_I6_n86, mult_42_I6_n85, mult_42_I6_n84, mult_42_I6_n83, 
      mult_42_I6_n82, mult_42_I6_n81, mult_42_I6_n80, mult_42_I6_n79, 
      mult_42_I6_n78, mult_42_I6_n77, mult_42_I6_n76, mult_42_I6_n75, 
      mult_42_I6_n74, mult_42_I6_n73, mult_42_I6_n72, mult_42_I6_n71, 
      mult_42_I6_n70, mult_42_I6_n69, mult_42_I6_n68, mult_42_I6_n67, 
      mult_42_I6_n66, mult_42_I6_n65, mult_42_I6_n64, mult_42_I6_n63, 
      mult_42_I6_n62, mult_42_I6_n61, mult_42_I6_n60, mult_42_I6_n59, 
      mult_42_I6_n58, mult_42_I6_n57, mult_42_I6_n56, mult_42_I6_n55, 
      mult_42_I6_n54, mult_42_I6_n53, mult_42_I6_n52, mult_42_I6_n51, 
      mult_42_I6_n50, mult_42_I6_n48, mult_42_I6_n47, mult_42_I6_n46, 
      mult_42_I6_n45, mult_42_I6_n44, mult_42_I6_n43, mult_42_I6_n42, 
      mult_42_I6_n41, mult_42_I6_n40, mult_42_I6_n39, mult_42_I6_n38, 
      mult_42_I6_n37, mult_42_I6_n35, mult_42_I6_n34, mult_42_I6_n33, 
      mult_42_I6_n32, mult_42_I6_n31, mult_42_I6_n30, mult_42_I6_n29, 
      mult_42_I6_n28, mult_42_I6_n27, mult_42_I6_n25, mult_42_I6_n24, 
      mult_42_I6_n23, mult_42_I6_n22, mult_42_I6_n21, mult_42_I6_n19, 
      mult_42_I6_n10, mult_42_I6_n9, mult_42_I6_n8, mult_42_I6_n7, 
      mult_42_I6_n6, mult_42_I6_n5, mult_42_I6_n4, mult_42_I6_n3, mult_42_I6_n2
      , mult_42_I6_n1, mult_42_I7_n402, mult_42_I7_n401, mult_42_I7_n400, 
      mult_42_I7_n399, mult_42_I7_n398, mult_42_I7_n397, mult_42_I7_n396, 
      mult_42_I7_n395, mult_42_I7_n394, mult_42_I7_n393, mult_42_I7_n392, 
      mult_42_I7_n391, mult_42_I7_n390, mult_42_I7_n389, mult_42_I7_n388, 
      mult_42_I7_n387, mult_42_I7_n386, mult_42_I7_n385, mult_42_I7_n384, 
      mult_42_I7_n383, mult_42_I7_n382, mult_42_I7_n381, mult_42_I7_n380, 
      mult_42_I7_n379, mult_42_I7_n378, mult_42_I7_n377, mult_42_I7_n376, 
      mult_42_I7_n375, mult_42_I7_n374, mult_42_I7_n373, mult_42_I7_n372, 
      mult_42_I7_n371, mult_42_I7_n370, mult_42_I7_n369, mult_42_I7_n368, 
      mult_42_I7_n367, mult_42_I7_n366, mult_42_I7_n365, mult_42_I7_n364, 
      mult_42_I7_n363, mult_42_I7_n362, mult_42_I7_n361, mult_42_I7_n360, 
      mult_42_I7_n359, mult_42_I7_n358, mult_42_I7_n357, mult_42_I7_n356, 
      mult_42_I7_n355, mult_42_I7_n354, mult_42_I7_n353, mult_42_I7_n352, 
      mult_42_I7_n351, mult_42_I7_n350, mult_42_I7_n349, mult_42_I7_n348, 
      mult_42_I7_n347, mult_42_I7_n346, mult_42_I7_n345, mult_42_I7_n344, 
      mult_42_I7_n343, mult_42_I7_n342, mult_42_I7_n341, mult_42_I7_n340, 
      mult_42_I7_n339, mult_42_I7_n338, mult_42_I7_n337, mult_42_I7_n336, 
      mult_42_I7_n335, mult_42_I7_n334, mult_42_I7_n333, mult_42_I7_n332, 
      mult_42_I7_n331, mult_42_I7_n330, mult_42_I7_n329, mult_42_I7_n328, 
      mult_42_I7_n327, mult_42_I7_n326, mult_42_I7_n325, mult_42_I7_n324, 
      mult_42_I7_n323, mult_42_I7_n322, mult_42_I7_n321, mult_42_I7_n320, 
      mult_42_I7_n319, mult_42_I7_n318, mult_42_I7_n317, mult_42_I7_n316, 
      mult_42_I7_n315, mult_42_I7_n314, mult_42_I7_n313, mult_42_I7_n312, 
      mult_42_I7_n311, mult_42_I7_n310, mult_42_I7_n309, mult_42_I7_n308, 
      mult_42_I7_n307, mult_42_I7_n306, mult_42_I7_n305, mult_42_I7_n304, 
      mult_42_I7_n303, mult_42_I7_n302, mult_42_I7_n301, mult_42_I7_n300, 
      mult_42_I7_n299, mult_42_I7_n298, mult_42_I7_n297, mult_42_I7_n296, 
      mult_42_I7_n295, mult_42_I7_n157, mult_42_I7_n156, mult_42_I7_n155, 
      mult_42_I7_n154, mult_42_I7_n153, mult_42_I7_n152, mult_42_I7_n151, 
      mult_42_I7_n148, mult_42_I7_n147, mult_42_I7_n146, mult_42_I7_n145, 
      mult_42_I7_n144, mult_42_I7_n143, mult_42_I7_n142, mult_42_I7_n140, 
      mult_42_I7_n139, mult_42_I7_n138, mult_42_I7_n137, mult_42_I7_n136, 
      mult_42_I7_n135, mult_42_I7_n134, mult_42_I7_n133, mult_42_I7_n132, 
      mult_42_I7_n131, mult_42_I7_n129, mult_42_I7_n128, mult_42_I7_n127, 
      mult_42_I7_n126, mult_42_I7_n124, mult_42_I7_n123, mult_42_I7_n122, 
      mult_42_I7_n121, mult_42_I7_n119, mult_42_I7_n118, mult_42_I7_n117, 
      mult_42_I7_n116, mult_42_I7_n115, mult_42_I7_n114, mult_42_I7_n113, 
      mult_42_I7_n112, mult_42_I7_n111, mult_42_I7_n107, mult_42_I7_n106, 
      mult_42_I7_n105, mult_42_I7_n90, mult_42_I7_n89, mult_42_I7_n88, 
      mult_42_I7_n87, mult_42_I7_n86, mult_42_I7_n85, mult_42_I7_n84, 
      mult_42_I7_n83, mult_42_I7_n82, mult_42_I7_n81, mult_42_I7_n80, 
      mult_42_I7_n79, mult_42_I7_n78, mult_42_I7_n77, mult_42_I7_n76, 
      mult_42_I7_n75, mult_42_I7_n74, mult_42_I7_n73, mult_42_I7_n72, 
      mult_42_I7_n71, mult_42_I7_n70, mult_42_I7_n69, mult_42_I7_n68, 
      mult_42_I7_n67, mult_42_I7_n66, mult_42_I7_n65, mult_42_I7_n64, 
      mult_42_I7_n63, mult_42_I7_n62, mult_42_I7_n61, mult_42_I7_n60, 
      mult_42_I7_n59, mult_42_I7_n58, mult_42_I7_n57, mult_42_I7_n56, 
      mult_42_I7_n55, mult_42_I7_n54, mult_42_I7_n53, mult_42_I7_n52, 
      mult_42_I7_n51, mult_42_I7_n50, mult_42_I7_n48, mult_42_I7_n47, 
      mult_42_I7_n46, mult_42_I7_n45, mult_42_I7_n44, mult_42_I7_n43, 
      mult_42_I7_n42, mult_42_I7_n41, mult_42_I7_n40, mult_42_I7_n39, 
      mult_42_I7_n38, mult_42_I7_n37, mult_42_I7_n35, mult_42_I7_n34, 
      mult_42_I7_n33, mult_42_I7_n32, mult_42_I7_n31, mult_42_I7_n30, 
      mult_42_I7_n29, mult_42_I7_n28, mult_42_I7_n27, mult_42_I7_n25, 
      mult_42_I7_n24, mult_42_I7_n23, mult_42_I7_n22, mult_42_I7_n21, 
      mult_42_I7_n19, mult_42_I7_n10, mult_42_I7_n9, mult_42_I7_n8, 
      mult_42_I7_n7, mult_42_I7_n6, mult_42_I7_n5, mult_42_I7_n4, mult_42_I7_n3
      , mult_42_I7_n2, mult_42_I7_n1, mult_42_I8_n402, mult_42_I8_n401, 
      mult_42_I8_n400, mult_42_I8_n399, mult_42_I8_n398, mult_42_I8_n397, 
      mult_42_I8_n396, mult_42_I8_n395, mult_42_I8_n394, mult_42_I8_n393, 
      mult_42_I8_n392, mult_42_I8_n391, mult_42_I8_n390, mult_42_I8_n389, 
      mult_42_I8_n388, mult_42_I8_n387, mult_42_I8_n386, mult_42_I8_n385, 
      mult_42_I8_n384, mult_42_I8_n383, mult_42_I8_n382, mult_42_I8_n381, 
      mult_42_I8_n380, mult_42_I8_n379, mult_42_I8_n378, mult_42_I8_n377, 
      mult_42_I8_n376, mult_42_I8_n375, mult_42_I8_n374, mult_42_I8_n373, 
      mult_42_I8_n372, mult_42_I8_n371, mult_42_I8_n370, mult_42_I8_n369, 
      mult_42_I8_n368, mult_42_I8_n367, mult_42_I8_n366, mult_42_I8_n365, 
      mult_42_I8_n364, mult_42_I8_n363, mult_42_I8_n362, mult_42_I8_n361, 
      mult_42_I8_n360, mult_42_I8_n359, mult_42_I8_n358, mult_42_I8_n357, 
      mult_42_I8_n356, mult_42_I8_n355, mult_42_I8_n354, mult_42_I8_n353, 
      mult_42_I8_n352, mult_42_I8_n351, mult_42_I8_n350, mult_42_I8_n349, 
      mult_42_I8_n348, mult_42_I8_n347, mult_42_I8_n346, mult_42_I8_n345, 
      mult_42_I8_n344, mult_42_I8_n343, mult_42_I8_n342, mult_42_I8_n341, 
      mult_42_I8_n340, mult_42_I8_n339, mult_42_I8_n338, mult_42_I8_n337, 
      mult_42_I8_n336, mult_42_I8_n335, mult_42_I8_n334, mult_42_I8_n333, 
      mult_42_I8_n332, mult_42_I8_n331, mult_42_I8_n330, mult_42_I8_n329, 
      mult_42_I8_n328, mult_42_I8_n327, mult_42_I8_n326, mult_42_I8_n325, 
      mult_42_I8_n324, mult_42_I8_n323, mult_42_I8_n322, mult_42_I8_n321, 
      mult_42_I8_n320, mult_42_I8_n319, mult_42_I8_n318, mult_42_I8_n317, 
      mult_42_I8_n316, mult_42_I8_n315, mult_42_I8_n314, mult_42_I8_n313, 
      mult_42_I8_n312, mult_42_I8_n311, mult_42_I8_n310, mult_42_I8_n309, 
      mult_42_I8_n308, mult_42_I8_n307, mult_42_I8_n306, mult_42_I8_n305, 
      mult_42_I8_n304, mult_42_I8_n303, mult_42_I8_n302, mult_42_I8_n301, 
      mult_42_I8_n300, mult_42_I8_n299, mult_42_I8_n298, mult_42_I8_n297, 
      mult_42_I8_n296, mult_42_I8_n295, mult_42_I8_n157, mult_42_I8_n156, 
      mult_42_I8_n155, mult_42_I8_n154, mult_42_I8_n153, mult_42_I8_n152, 
      mult_42_I8_n151, mult_42_I8_n148, mult_42_I8_n147, mult_42_I8_n146, 
      mult_42_I8_n145, mult_42_I8_n144, mult_42_I8_n143, mult_42_I8_n142, 
      mult_42_I8_n140, mult_42_I8_n139, mult_42_I8_n138, mult_42_I8_n137, 
      mult_42_I8_n136, mult_42_I8_n135, mult_42_I8_n134, mult_42_I8_n133, 
      mult_42_I8_n132, mult_42_I8_n131, mult_42_I8_n129, mult_42_I8_n128, 
      mult_42_I8_n127, mult_42_I8_n126, mult_42_I8_n124, mult_42_I8_n123, 
      mult_42_I8_n122, mult_42_I8_n121, mult_42_I8_n119, mult_42_I8_n118, 
      mult_42_I8_n117, mult_42_I8_n116, mult_42_I8_n115, mult_42_I8_n114, 
      mult_42_I8_n113, mult_42_I8_n112, mult_42_I8_n111, mult_42_I8_n107, 
      mult_42_I8_n106, mult_42_I8_n105, mult_42_I8_n90, mult_42_I8_n89, 
      mult_42_I8_n88, mult_42_I8_n87, mult_42_I8_n86, mult_42_I8_n85, 
      mult_42_I8_n84, mult_42_I8_n83, mult_42_I8_n82, mult_42_I8_n81, 
      mult_42_I8_n80, mult_42_I8_n79, mult_42_I8_n78, mult_42_I8_n77, 
      mult_42_I8_n76, mult_42_I8_n75, mult_42_I8_n74, mult_42_I8_n73, 
      mult_42_I8_n72, mult_42_I8_n71, mult_42_I8_n70, mult_42_I8_n69, 
      mult_42_I8_n68, mult_42_I8_n67, mult_42_I8_n66, mult_42_I8_n65, 
      mult_42_I8_n64, mult_42_I8_n63, mult_42_I8_n62, mult_42_I8_n61, 
      mult_42_I8_n60, mult_42_I8_n59, mult_42_I8_n58, mult_42_I8_n57, 
      mult_42_I8_n56, mult_42_I8_n55, mult_42_I8_n54, mult_42_I8_n53, 
      mult_42_I8_n52, mult_42_I8_n51, mult_42_I8_n50, mult_42_I8_n48, 
      mult_42_I8_n47, mult_42_I8_n46, mult_42_I8_n45, mult_42_I8_n44, 
      mult_42_I8_n43, mult_42_I8_n42, mult_42_I8_n41, mult_42_I8_n40, 
      mult_42_I8_n39, mult_42_I8_n38, mult_42_I8_n37, mult_42_I8_n35, 
      mult_42_I8_n34, mult_42_I8_n33, mult_42_I8_n32, mult_42_I8_n31, 
      mult_42_I8_n30, mult_42_I8_n29, mult_42_I8_n28, mult_42_I8_n27, 
      mult_42_I8_n25, mult_42_I8_n24, mult_42_I8_n23, mult_42_I8_n22, 
      mult_42_I8_n21, mult_42_I8_n19, mult_42_I8_n10, mult_42_I8_n9, 
      mult_42_I8_n8, mult_42_I8_n7, mult_42_I8_n6, mult_42_I8_n5, mult_42_I8_n4
      , mult_42_I8_n3, mult_42_I8_n2, mult_42_I8_n1, mult_42_I9_n402, 
      mult_42_I9_n401, mult_42_I9_n400, mult_42_I9_n399, mult_42_I9_n398, 
      mult_42_I9_n397, mult_42_I9_n396, mult_42_I9_n395, mult_42_I9_n394, 
      mult_42_I9_n393, mult_42_I9_n392, mult_42_I9_n391, mult_42_I9_n390, 
      mult_42_I9_n389, mult_42_I9_n388, mult_42_I9_n387, mult_42_I9_n386, 
      mult_42_I9_n385, mult_42_I9_n384, mult_42_I9_n383, mult_42_I9_n382, 
      mult_42_I9_n381, mult_42_I9_n380, mult_42_I9_n379, mult_42_I9_n378, 
      mult_42_I9_n377, mult_42_I9_n376, mult_42_I9_n375, mult_42_I9_n374, 
      mult_42_I9_n373, mult_42_I9_n372, mult_42_I9_n371, mult_42_I9_n370, 
      mult_42_I9_n369, mult_42_I9_n368, mult_42_I9_n367, mult_42_I9_n366, 
      mult_42_I9_n365, mult_42_I9_n364, mult_42_I9_n363, mult_42_I9_n362, 
      mult_42_I9_n361, mult_42_I9_n360, mult_42_I9_n359, mult_42_I9_n358, 
      mult_42_I9_n357, mult_42_I9_n356, mult_42_I9_n355, mult_42_I9_n354, 
      mult_42_I9_n353, mult_42_I9_n352, mult_42_I9_n351, mult_42_I9_n350, 
      mult_42_I9_n349, mult_42_I9_n348, mult_42_I9_n347, mult_42_I9_n346, 
      mult_42_I9_n345, mult_42_I9_n344, mult_42_I9_n343, mult_42_I9_n342, 
      mult_42_I9_n341, mult_42_I9_n340, mult_42_I9_n339, mult_42_I9_n338, 
      mult_42_I9_n337, mult_42_I9_n336, mult_42_I9_n335, mult_42_I9_n334, 
      mult_42_I9_n333, mult_42_I9_n332, mult_42_I9_n331, mult_42_I9_n330, 
      mult_42_I9_n329, mult_42_I9_n328, mult_42_I9_n327, mult_42_I9_n326, 
      mult_42_I9_n325, mult_42_I9_n324, mult_42_I9_n323, mult_42_I9_n322, 
      mult_42_I9_n321, mult_42_I9_n320, mult_42_I9_n319, mult_42_I9_n318, 
      mult_42_I9_n317, mult_42_I9_n316, mult_42_I9_n315, mult_42_I9_n314, 
      mult_42_I9_n313, mult_42_I9_n312, mult_42_I9_n311, mult_42_I9_n310, 
      mult_42_I9_n309, mult_42_I9_n308, mult_42_I9_n307, mult_42_I9_n306, 
      mult_42_I9_n305, mult_42_I9_n304, mult_42_I9_n303, mult_42_I9_n302, 
      mult_42_I9_n301, mult_42_I9_n300, mult_42_I9_n299, mult_42_I9_n298, 
      mult_42_I9_n297, mult_42_I9_n296, mult_42_I9_n295, mult_42_I9_n157, 
      mult_42_I9_n156, mult_42_I9_n155, mult_42_I9_n154, mult_42_I9_n153, 
      mult_42_I9_n152, mult_42_I9_n151, mult_42_I9_n148, mult_42_I9_n147, 
      mult_42_I9_n146, mult_42_I9_n145, mult_42_I9_n144, mult_42_I9_n143, 
      mult_42_I9_n142, mult_42_I9_n140, mult_42_I9_n139, mult_42_I9_n138, 
      mult_42_I9_n137, mult_42_I9_n136, mult_42_I9_n135, mult_42_I9_n134, 
      mult_42_I9_n133, mult_42_I9_n132, mult_42_I9_n131, mult_42_I9_n129, 
      mult_42_I9_n128, mult_42_I9_n127, mult_42_I9_n126, mult_42_I9_n124, 
      mult_42_I9_n123, mult_42_I9_n122, mult_42_I9_n121, mult_42_I9_n119, 
      mult_42_I9_n118, mult_42_I9_n117, mult_42_I9_n116, mult_42_I9_n115, 
      mult_42_I9_n114, mult_42_I9_n113, mult_42_I9_n112, mult_42_I9_n111, 
      mult_42_I9_n107, mult_42_I9_n106, mult_42_I9_n105, mult_42_I9_n90, 
      mult_42_I9_n89, mult_42_I9_n88, mult_42_I9_n87, mult_42_I9_n86, 
      mult_42_I9_n85, mult_42_I9_n84, mult_42_I9_n83, mult_42_I9_n82, 
      mult_42_I9_n81, mult_42_I9_n80, mult_42_I9_n79, mult_42_I9_n78, 
      mult_42_I9_n77, mult_42_I9_n76, mult_42_I9_n75, mult_42_I9_n74, 
      mult_42_I9_n73, mult_42_I9_n72, mult_42_I9_n71, mult_42_I9_n70, 
      mult_42_I9_n69, mult_42_I9_n68, mult_42_I9_n67, mult_42_I9_n66, 
      mult_42_I9_n65, mult_42_I9_n64, mult_42_I9_n63, mult_42_I9_n62, 
      mult_42_I9_n61, mult_42_I9_n60, mult_42_I9_n59, mult_42_I9_n58, 
      mult_42_I9_n57, mult_42_I9_n56, mult_42_I9_n55, mult_42_I9_n54, 
      mult_42_I9_n53, mult_42_I9_n52, mult_42_I9_n51, mult_42_I9_n50, 
      mult_42_I9_n48, mult_42_I9_n47, mult_42_I9_n46, mult_42_I9_n45, 
      mult_42_I9_n44, mult_42_I9_n43, mult_42_I9_n42, mult_42_I9_n41, 
      mult_42_I9_n40, mult_42_I9_n39, mult_42_I9_n38, mult_42_I9_n37, 
      mult_42_I9_n35, mult_42_I9_n34, mult_42_I9_n33, mult_42_I9_n32, 
      mult_42_I9_n31, mult_42_I9_n30, mult_42_I9_n29, mult_42_I9_n28, 
      mult_42_I9_n27, mult_42_I9_n25, mult_42_I9_n24, mult_42_I9_n23, 
      mult_42_I9_n22, mult_42_I9_n21, mult_42_I9_n19, mult_42_I9_n10, 
      mult_42_I9_n9, mult_42_I9_n8, mult_42_I9_n7, mult_42_I9_n6, mult_42_I9_n5
      , mult_42_I9_n4, mult_42_I9_n3, mult_42_I9_n2, mult_42_I9_n1, 
      mult_42_I10_n402, mult_42_I10_n401, mult_42_I10_n400, mult_42_I10_n399, 
      mult_42_I10_n398, mult_42_I10_n397, mult_42_I10_n396, mult_42_I10_n395, 
      mult_42_I10_n394, mult_42_I10_n393, mult_42_I10_n392, mult_42_I10_n391, 
      mult_42_I10_n390, mult_42_I10_n389, mult_42_I10_n388, mult_42_I10_n387, 
      mult_42_I10_n386, mult_42_I10_n385, mult_42_I10_n384, mult_42_I10_n383, 
      mult_42_I10_n382, mult_42_I10_n381, mult_42_I10_n380, mult_42_I10_n379, 
      mult_42_I10_n378, mult_42_I10_n377, mult_42_I10_n376, mult_42_I10_n375, 
      mult_42_I10_n374, mult_42_I10_n373, mult_42_I10_n372, mult_42_I10_n371, 
      mult_42_I10_n370, mult_42_I10_n369, mult_42_I10_n368, mult_42_I10_n367, 
      mult_42_I10_n366, mult_42_I10_n365, mult_42_I10_n364, mult_42_I10_n363, 
      mult_42_I10_n362, mult_42_I10_n361, mult_42_I10_n360, mult_42_I10_n359, 
      mult_42_I10_n358, mult_42_I10_n357, mult_42_I10_n356, mult_42_I10_n355, 
      mult_42_I10_n354, mult_42_I10_n353, mult_42_I10_n352, mult_42_I10_n351, 
      mult_42_I10_n350, mult_42_I10_n349, mult_42_I10_n348, mult_42_I10_n347, 
      mult_42_I10_n346, mult_42_I10_n345, mult_42_I10_n344, mult_42_I10_n343, 
      mult_42_I10_n342, mult_42_I10_n341, mult_42_I10_n340, mult_42_I10_n339, 
      mult_42_I10_n338, mult_42_I10_n337, mult_42_I10_n336, mult_42_I10_n335, 
      mult_42_I10_n334, mult_42_I10_n333, mult_42_I10_n332, mult_42_I10_n331, 
      mult_42_I10_n330, mult_42_I10_n329, mult_42_I10_n328, mult_42_I10_n327, 
      mult_42_I10_n326, mult_42_I10_n325, mult_42_I10_n324, mult_42_I10_n323, 
      mult_42_I10_n322, mult_42_I10_n321, mult_42_I10_n320, mult_42_I10_n319, 
      mult_42_I10_n318, mult_42_I10_n317, mult_42_I10_n316, mult_42_I10_n315, 
      mult_42_I10_n314, mult_42_I10_n313, mult_42_I10_n312, mult_42_I10_n311, 
      mult_42_I10_n310, mult_42_I10_n309, mult_42_I10_n308, mult_42_I10_n307, 
      mult_42_I10_n306, mult_42_I10_n305, mult_42_I10_n304, mult_42_I10_n303, 
      mult_42_I10_n302, mult_42_I10_n301, mult_42_I10_n300, mult_42_I10_n299, 
      mult_42_I10_n298, mult_42_I10_n297, mult_42_I10_n296, mult_42_I10_n295, 
      mult_42_I10_n157, mult_42_I10_n156, mult_42_I10_n155, mult_42_I10_n154, 
      mult_42_I10_n153, mult_42_I10_n152, mult_42_I10_n151, mult_42_I10_n148, 
      mult_42_I10_n147, mult_42_I10_n146, mult_42_I10_n145, mult_42_I10_n144, 
      mult_42_I10_n143, mult_42_I10_n142, mult_42_I10_n140, mult_42_I10_n139, 
      mult_42_I10_n138, mult_42_I10_n137, mult_42_I10_n136, mult_42_I10_n135, 
      mult_42_I10_n134, mult_42_I10_n133, mult_42_I10_n132, mult_42_I10_n131, 
      mult_42_I10_n129, mult_42_I10_n128, mult_42_I10_n127, mult_42_I10_n126, 
      mult_42_I10_n124, mult_42_I10_n123, mult_42_I10_n122, mult_42_I10_n121, 
      mult_42_I10_n119, mult_42_I10_n118, mult_42_I10_n117, mult_42_I10_n116, 
      mult_42_I10_n115, mult_42_I10_n114, mult_42_I10_n113, mult_42_I10_n112, 
      mult_42_I10_n111, mult_42_I10_n107, mult_42_I10_n106, mult_42_I10_n105, 
      mult_42_I10_n90, mult_42_I10_n89, mult_42_I10_n88, mult_42_I10_n87, 
      mult_42_I10_n86, mult_42_I10_n85, mult_42_I10_n84, mult_42_I10_n83, 
      mult_42_I10_n82, mult_42_I10_n81, mult_42_I10_n80, mult_42_I10_n79, 
      mult_42_I10_n78, mult_42_I10_n77, mult_42_I10_n76, mult_42_I10_n75, 
      mult_42_I10_n74, mult_42_I10_n73, mult_42_I10_n72, mult_42_I10_n71, 
      mult_42_I10_n70, mult_42_I10_n69, mult_42_I10_n68, mult_42_I10_n67, 
      mult_42_I10_n66, mult_42_I10_n65, mult_42_I10_n64, mult_42_I10_n63, 
      mult_42_I10_n62, mult_42_I10_n61, mult_42_I10_n60, mult_42_I10_n59, 
      mult_42_I10_n58, mult_42_I10_n57, mult_42_I10_n56, mult_42_I10_n55, 
      mult_42_I10_n54, mult_42_I10_n53, mult_42_I10_n52, mult_42_I10_n51, 
      mult_42_I10_n50, mult_42_I10_n48, mult_42_I10_n47, mult_42_I10_n46, 
      mult_42_I10_n45, mult_42_I10_n44, mult_42_I10_n43, mult_42_I10_n42, 
      mult_42_I10_n41, mult_42_I10_n40, mult_42_I10_n39, mult_42_I10_n38, 
      mult_42_I10_n37, mult_42_I10_n35, mult_42_I10_n34, mult_42_I10_n33, 
      mult_42_I10_n32, mult_42_I10_n31, mult_42_I10_n30, mult_42_I10_n29, 
      mult_42_I10_n28, mult_42_I10_n27, mult_42_I10_n25, mult_42_I10_n24, 
      mult_42_I10_n23, mult_42_I10_n22, mult_42_I10_n21, mult_42_I10_n19, 
      mult_42_I10_n10, mult_42_I10_n9, mult_42_I10_n8, mult_42_I10_n7, 
      mult_42_I10_n6, mult_42_I10_n5, mult_42_I10_n4, mult_42_I10_n3, 
      mult_42_I10_n2, mult_42_I10_n1, mult_42_I11_n402, mult_42_I11_n401, 
      mult_42_I11_n400, mult_42_I11_n399, mult_42_I11_n398, mult_42_I11_n397, 
      mult_42_I11_n396, mult_42_I11_n395, mult_42_I11_n394, mult_42_I11_n393, 
      mult_42_I11_n392, mult_42_I11_n391, mult_42_I11_n390, mult_42_I11_n389, 
      mult_42_I11_n388, mult_42_I11_n387, mult_42_I11_n386, mult_42_I11_n385, 
      mult_42_I11_n384, mult_42_I11_n383, mult_42_I11_n382, mult_42_I11_n381, 
      mult_42_I11_n380, mult_42_I11_n379, mult_42_I11_n378, mult_42_I11_n377, 
      mult_42_I11_n376, mult_42_I11_n375, mult_42_I11_n374, mult_42_I11_n373, 
      mult_42_I11_n372, mult_42_I11_n371, mult_42_I11_n370, mult_42_I11_n369, 
      mult_42_I11_n368, mult_42_I11_n367, mult_42_I11_n366, mult_42_I11_n365, 
      mult_42_I11_n364, mult_42_I11_n363, mult_42_I11_n362, mult_42_I11_n361, 
      mult_42_I11_n360, mult_42_I11_n359, mult_42_I11_n358, mult_42_I11_n357, 
      mult_42_I11_n356, mult_42_I11_n355, mult_42_I11_n354, mult_42_I11_n353, 
      mult_42_I11_n352, mult_42_I11_n351, mult_42_I11_n350, mult_42_I11_n349, 
      mult_42_I11_n348, mult_42_I11_n347, mult_42_I11_n346, mult_42_I11_n345, 
      mult_42_I11_n344, mult_42_I11_n343, mult_42_I11_n342, mult_42_I11_n341, 
      mult_42_I11_n340, mult_42_I11_n339, mult_42_I11_n338, mult_42_I11_n337, 
      mult_42_I11_n336, mult_42_I11_n335, mult_42_I11_n334, mult_42_I11_n333, 
      mult_42_I11_n332, mult_42_I11_n331, mult_42_I11_n330, mult_42_I11_n329, 
      mult_42_I11_n328, mult_42_I11_n327, mult_42_I11_n326, mult_42_I11_n325, 
      mult_42_I11_n324, mult_42_I11_n323, mult_42_I11_n322, mult_42_I11_n321, 
      mult_42_I11_n320, mult_42_I11_n319, mult_42_I11_n318, mult_42_I11_n317, 
      mult_42_I11_n316, mult_42_I11_n315, mult_42_I11_n314, mult_42_I11_n313, 
      mult_42_I11_n312, mult_42_I11_n311, mult_42_I11_n310, mult_42_I11_n309, 
      mult_42_I11_n308, mult_42_I11_n307, mult_42_I11_n306, mult_42_I11_n305, 
      mult_42_I11_n304, mult_42_I11_n303, mult_42_I11_n302, mult_42_I11_n301, 
      mult_42_I11_n300, mult_42_I11_n299, mult_42_I11_n298, mult_42_I11_n297, 
      mult_42_I11_n296, mult_42_I11_n295, mult_42_I11_n157, mult_42_I11_n156, 
      mult_42_I11_n155, mult_42_I11_n154, mult_42_I11_n153, mult_42_I11_n152, 
      mult_42_I11_n151, mult_42_I11_n148, mult_42_I11_n147, mult_42_I11_n146, 
      mult_42_I11_n145, mult_42_I11_n144, mult_42_I11_n143, mult_42_I11_n142, 
      mult_42_I11_n140, mult_42_I11_n139, mult_42_I11_n138, mult_42_I11_n137, 
      mult_42_I11_n136, mult_42_I11_n135, mult_42_I11_n134, mult_42_I11_n133, 
      mult_42_I11_n132, mult_42_I11_n131, mult_42_I11_n129, mult_42_I11_n128, 
      mult_42_I11_n127, mult_42_I11_n126, mult_42_I11_n124, mult_42_I11_n123, 
      mult_42_I11_n122, mult_42_I11_n121, mult_42_I11_n119, mult_42_I11_n118, 
      mult_42_I11_n117, mult_42_I11_n116, mult_42_I11_n115, mult_42_I11_n114, 
      mult_42_I11_n113, mult_42_I11_n112, mult_42_I11_n111, mult_42_I11_n107, 
      mult_42_I11_n106, mult_42_I11_n105, mult_42_I11_n90, mult_42_I11_n89, 
      mult_42_I11_n88, mult_42_I11_n87, mult_42_I11_n86, mult_42_I11_n85, 
      mult_42_I11_n84, mult_42_I11_n83, mult_42_I11_n82, mult_42_I11_n81, 
      mult_42_I11_n80, mult_42_I11_n79, mult_42_I11_n78, mult_42_I11_n77, 
      mult_42_I11_n76, mult_42_I11_n75, mult_42_I11_n74, mult_42_I11_n73, 
      mult_42_I11_n72, mult_42_I11_n71, mult_42_I11_n70, mult_42_I11_n69, 
      mult_42_I11_n68, mult_42_I11_n67, mult_42_I11_n66, mult_42_I11_n65, 
      mult_42_I11_n64, mult_42_I11_n63, mult_42_I11_n62, mult_42_I11_n61, 
      mult_42_I11_n60, mult_42_I11_n59, mult_42_I11_n58, mult_42_I11_n57, 
      mult_42_I11_n56, mult_42_I11_n55, mult_42_I11_n54, mult_42_I11_n53, 
      mult_42_I11_n52, mult_42_I11_n51, mult_42_I11_n50, mult_42_I11_n48, 
      mult_42_I11_n47, mult_42_I11_n46, mult_42_I11_n45, mult_42_I11_n44, 
      mult_42_I11_n43, mult_42_I11_n42, mult_42_I11_n41, mult_42_I11_n40, 
      mult_42_I11_n39, mult_42_I11_n38, mult_42_I11_n37, mult_42_I11_n35, 
      mult_42_I11_n34, mult_42_I11_n33, mult_42_I11_n32, mult_42_I11_n31, 
      mult_42_I11_n30, mult_42_I11_n29, mult_42_I11_n28, mult_42_I11_n27, 
      mult_42_I11_n25, mult_42_I11_n24, mult_42_I11_n23, mult_42_I11_n22, 
      mult_42_I11_n21, mult_42_I11_n19, mult_42_I11_n10, mult_42_I11_n9, 
      mult_42_I11_n8, mult_42_I11_n7, mult_42_I11_n6, mult_42_I11_n5, 
      mult_42_I11_n4, mult_42_I11_n3, mult_42_I11_n2, mult_42_I11_n1, 
      add_6_root_add_0_root_add_44_I11_n_1112, 
      add_6_root_add_0_root_add_44_I11_n1, 
      add_6_root_add_0_root_add_44_I11_carry_2_port, 
      add_6_root_add_0_root_add_44_I11_carry_3_port, 
      add_6_root_add_0_root_add_44_I11_carry_4_port, 
      add_6_root_add_0_root_add_44_I11_carry_5_port, 
      add_6_root_add_0_root_add_44_I11_carry_6_port, 
      add_6_root_add_0_root_add_44_I11_carry_7_port, 
      add_6_root_add_0_root_add_44_I11_carry_8_port, 
      add_6_root_add_0_root_add_44_I11_carry_9_port, 
      add_8_root_add_0_root_add_44_I11_n_1115, 
      add_8_root_add_0_root_add_44_I11_n1, 
      add_8_root_add_0_root_add_44_I11_carry_2_port, 
      add_8_root_add_0_root_add_44_I11_carry_3_port, 
      add_8_root_add_0_root_add_44_I11_carry_4_port, 
      add_8_root_add_0_root_add_44_I11_carry_5_port, 
      add_8_root_add_0_root_add_44_I11_carry_6_port, 
      add_8_root_add_0_root_add_44_I11_carry_7_port, 
      add_8_root_add_0_root_add_44_I11_carry_8_port, 
      add_8_root_add_0_root_add_44_I11_carry_9_port, 
      add_9_root_add_0_root_add_44_I11_n_1118, 
      add_9_root_add_0_root_add_44_I11_n1, 
      add_9_root_add_0_root_add_44_I11_carry_2_port, 
      add_9_root_add_0_root_add_44_I11_carry_3_port, 
      add_9_root_add_0_root_add_44_I11_carry_4_port, 
      add_9_root_add_0_root_add_44_I11_carry_5_port, 
      add_9_root_add_0_root_add_44_I11_carry_6_port, 
      add_9_root_add_0_root_add_44_I11_carry_7_port, 
      add_9_root_add_0_root_add_44_I11_carry_8_port, 
      add_9_root_add_0_root_add_44_I11_carry_9_port, 
      add_7_root_add_0_root_add_44_I11_n_1121, 
      add_7_root_add_0_root_add_44_I11_n1, 
      add_7_root_add_0_root_add_44_I11_carry_2_port, 
      add_7_root_add_0_root_add_44_I11_carry_3_port, 
      add_7_root_add_0_root_add_44_I11_carry_4_port, 
      add_7_root_add_0_root_add_44_I11_carry_5_port, 
      add_7_root_add_0_root_add_44_I11_carry_6_port, 
      add_7_root_add_0_root_add_44_I11_carry_7_port, 
      add_7_root_add_0_root_add_44_I11_carry_8_port, 
      add_7_root_add_0_root_add_44_I11_carry_9_port, 
      add_2_root_add_0_root_add_44_I11_n_1124, 
      add_2_root_add_0_root_add_44_I11_n1, 
      add_2_root_add_0_root_add_44_I11_carry_2_port, 
      add_2_root_add_0_root_add_44_I11_carry_3_port, 
      add_2_root_add_0_root_add_44_I11_carry_4_port, 
      add_2_root_add_0_root_add_44_I11_carry_5_port, 
      add_2_root_add_0_root_add_44_I11_carry_6_port, 
      add_2_root_add_0_root_add_44_I11_carry_7_port, 
      add_2_root_add_0_root_add_44_I11_carry_8_port, 
      add_2_root_add_0_root_add_44_I11_carry_9_port, 
      add_3_root_add_0_root_add_44_I11_n_1127, 
      add_3_root_add_0_root_add_44_I11_n1, 
      add_3_root_add_0_root_add_44_I11_carry_2_port, 
      add_3_root_add_0_root_add_44_I11_carry_3_port, 
      add_3_root_add_0_root_add_44_I11_carry_4_port, 
      add_3_root_add_0_root_add_44_I11_carry_5_port, 
      add_3_root_add_0_root_add_44_I11_carry_6_port, 
      add_3_root_add_0_root_add_44_I11_carry_7_port, 
      add_3_root_add_0_root_add_44_I11_carry_8_port, 
      add_3_root_add_0_root_add_44_I11_carry_9_port, 
      add_5_root_add_0_root_add_44_I11_n_1130, 
      add_5_root_add_0_root_add_44_I11_n1, 
      add_5_root_add_0_root_add_44_I11_carry_2_port, 
      add_5_root_add_0_root_add_44_I11_carry_3_port, 
      add_5_root_add_0_root_add_44_I11_carry_4_port, 
      add_5_root_add_0_root_add_44_I11_carry_5_port, 
      add_5_root_add_0_root_add_44_I11_carry_6_port, 
      add_5_root_add_0_root_add_44_I11_carry_7_port, 
      add_5_root_add_0_root_add_44_I11_carry_8_port, 
      add_5_root_add_0_root_add_44_I11_carry_9_port, 
      add_4_root_add_0_root_add_44_I11_n_1133, 
      add_4_root_add_0_root_add_44_I11_n1, 
      add_4_root_add_0_root_add_44_I11_carry_2_port, 
      add_4_root_add_0_root_add_44_I11_carry_3_port, 
      add_4_root_add_0_root_add_44_I11_carry_4_port, 
      add_4_root_add_0_root_add_44_I11_carry_5_port, 
      add_4_root_add_0_root_add_44_I11_carry_6_port, 
      add_4_root_add_0_root_add_44_I11_carry_7_port, 
      add_4_root_add_0_root_add_44_I11_carry_8_port, 
      add_4_root_add_0_root_add_44_I11_carry_9_port, 
      add_1_root_add_0_root_add_44_I11_n_1136, 
      add_1_root_add_0_root_add_44_I11_n1, 
      add_1_root_add_0_root_add_44_I11_carry_2_port, 
      add_1_root_add_0_root_add_44_I11_carry_3_port, 
      add_1_root_add_0_root_add_44_I11_carry_4_port, 
      add_1_root_add_0_root_add_44_I11_carry_5_port, 
      add_1_root_add_0_root_add_44_I11_carry_6_port, 
      add_1_root_add_0_root_add_44_I11_carry_7_port, 
      add_1_root_add_0_root_add_44_I11_carry_8_port, 
      add_1_root_add_0_root_add_44_I11_carry_9_port, 
      add_0_root_add_0_root_add_44_I11_n_1139, 
      add_0_root_add_0_root_add_44_I11_n2, 
      add_0_root_add_0_root_add_44_I11_carry_2_port, 
      add_0_root_add_0_root_add_44_I11_carry_3_port, 
      add_0_root_add_0_root_add_44_I11_carry_4_port, 
      add_0_root_add_0_root_add_44_I11_carry_5_port, 
      add_0_root_add_0_root_add_44_I11_carry_6_port, 
      add_0_root_add_0_root_add_44_I11_carry_7_port, 
      add_0_root_add_0_root_add_44_I11_carry_8_port, 
      add_0_root_add_0_root_add_44_I11_carry_9_port : std_logic;

begin
   
   DOUT_reg_9_inst : DFF_X1 port map( D => n287, CK => clk, Q => DOUT(9), QN =>
                           n166);
   DOUT_reg_8_inst : DFF_X1 port map( D => n286, CK => clk, Q => DOUT(8), QN =>
                           n165);
   DOUT_reg_7_inst : DFF_X1 port map( D => n285, CK => clk, Q => DOUT(7), QN =>
                           n164);
   DOUT_reg_6_inst : DFF_X1 port map( D => n284, CK => clk, Q => DOUT(6), QN =>
                           n163);
   DOUT_reg_5_inst : DFF_X1 port map( D => n283, CK => clk, Q => DOUT(5), QN =>
                           n162);
   DOUT_reg_4_inst : DFF_X1 port map( D => n282, CK => clk, Q => DOUT(4), QN =>
                           n161);
   DOUT_reg_3_inst : DFF_X1 port map( D => n281, CK => clk, Q => DOUT(3), QN =>
                           n160);
   DOUT_reg_2_inst : DFF_X1 port map( D => n280, CK => clk, Q => DOUT(2), QN =>
                           n159);
   DOUT_reg_1_inst : DFF_X1 port map( D => n279, CK => clk, Q => DOUT(1), QN =>
                           n158);
   DOUT_reg_0_inst : DFF_X1 port map( D => n278, CK => clk, Q => DOUT(0), QN =>
                           n157);
   x_vector_reg_0_9_inst : DFF_X1 port map( D => n277, CK => clk, Q => 
                           x_vector_9_port, QN => n364);
   x_vector_reg_1_9_inst : DFF_X1 port map( D => n276, CK => clk, Q => 
                           x_vector_19_port, QN => n312);
   x_vector_reg_2_9_inst : DFF_X1 port map( D => n275, CK => clk, Q => 
                           x_vector_29_port, QN => n363);
   x_vector_reg_3_9_inst : DFF_X1 port map( D => n274, CK => clk, Q => 
                           x_vector_39_port, QN => n311);
   x_vector_reg_4_9_inst : DFF_X1 port map( D => n273, CK => clk, Q => 
                           x_vector_49_port, QN => n362);
   x_vector_reg_5_9_inst : DFF_X1 port map( D => n272, CK => clk, Q => 
                           x_vector_59_port, QN => n310);
   x_vector_reg_6_9_inst : DFF_X1 port map( D => n271, CK => clk, Q => 
                           x_vector_69_port, QN => n361);
   x_vector_reg_7_9_inst : DFF_X1 port map( D => n270, CK => clk, Q => 
                           x_vector_79_port, QN => n309);
   x_vector_reg_8_9_inst : DFF_X1 port map( D => n269, CK => clk, Q => 
                           x_vector_89_port, QN => n360);
   x_vector_reg_9_9_inst : DFF_X1 port map( D => n268, CK => clk, Q => 
                           x_vector_99_port, QN => n313);
   x_vector_reg_10_9_inst : DFF_X1 port map( D => n267, CK => clk, Q => 
                           x_vector_109_port, QN => n392);
   x_vector_reg_0_8_inst : DFF_X1 port map( D => n266, CK => clk, Q => 
                           x_vector_8_port, QN => n379);
   x_vector_reg_1_8_inst : DFF_X1 port map( D => n265, CK => clk, Q => 
                           x_vector_18_port, QN => n325);
   x_vector_reg_2_8_inst : DFF_X1 port map( D => n264, CK => clk, Q => 
                           x_vector_28_port, QN => n376);
   x_vector_reg_3_8_inst : DFF_X1 port map( D => n263, CK => clk, Q => 
                           x_vector_38_port, QN => n324);
   x_vector_reg_4_8_inst : DFF_X1 port map( D => n262, CK => clk, Q => 
                           x_vector_48_port, QN => n375);
   x_vector_reg_5_8_inst : DFF_X1 port map( D => n261, CK => clk, Q => 
                           x_vector_58_port, QN => n323);
   x_vector_reg_6_8_inst : DFF_X1 port map( D => n260, CK => clk, Q => 
                           x_vector_68_port, QN => n374);
   x_vector_reg_7_8_inst : DFF_X1 port map( D => n259, CK => clk, Q => 
                           x_vector_78_port, QN => n322);
   x_vector_reg_8_8_inst : DFF_X1 port map( D => n258, CK => clk, Q => 
                           x_vector_88_port, QN => n373);
   x_vector_reg_9_8_inst : DFF_X1 port map( D => n257, CK => clk, Q => 
                           x_vector_98_port, QN => n327);
   x_vector_reg_10_8_inst : DFF_X1 port map( D => n256, CK => clk, Q => 
                           x_vector_108_port, QN => n395);
   x_vector_reg_0_7_inst : DFF_X1 port map( D => n255, CK => clk, Q => 
                           x_vector_7_port, QN => n359);
   x_vector_reg_1_7_inst : DFF_X1 port map( D => n254, CK => clk, Q => 
                           x_vector_17_port, QN => n305);
   x_vector_reg_2_7_inst : DFF_X1 port map( D => n253, CK => clk, Q => 
                           x_vector_27_port, QN => n357);
   x_vector_reg_3_7_inst : DFF_X1 port map( D => n252, CK => clk, Q => 
                           x_vector_37_port, QN => n304);
   x_vector_reg_4_7_inst : DFF_X1 port map( D => n251, CK => clk, Q => 
                           x_vector_47_port, QN => n356);
   x_vector_reg_5_7_inst : DFF_X1 port map( D => n250, CK => clk, Q => 
                           x_vector_57_port, QN => n303);
   x_vector_reg_6_7_inst : DFF_X1 port map( D => n249, CK => clk, Q => 
                           x_vector_67_port, QN => n355);
   x_vector_reg_7_7_inst : DFF_X1 port map( D => n248, CK => clk, Q => 
                           x_vector_77_port, QN => n302);
   x_vector_reg_8_7_inst : DFF_X1 port map( D => n247, CK => clk, Q => 
                           x_vector_87_port, QN => n354);
   x_vector_reg_9_7_inst : DFF_X1 port map( D => n246, CK => clk, Q => 
                           x_vector_97_port, QN => n307);
   x_vector_reg_10_7_inst : DFF_X1 port map( D => n245, CK => clk, Q => 
                           x_vector_107_port, QN => n391);
   x_vector_reg_0_6_inst : DFF_X1 port map( D => n244, CK => clk, Q => 
                           x_vector_6_port, QN => n378);
   x_vector_reg_1_6_inst : DFF_X1 port map( D => n243, CK => clk, Q => 
                           x_vector_16_port, QN => n321);
   x_vector_reg_2_6_inst : DFF_X1 port map( D => n242, CK => clk, Q => 
                           x_vector_26_port, QN => n367);
   x_vector_reg_3_6_inst : DFF_X1 port map( D => n241, CK => clk, Q => 
                           x_vector_36_port, QN => n316);
   x_vector_reg_4_6_inst : DFF_X1 port map( D => n240, CK => clk, Q => 
                           x_vector_46_port, QN => n366);
   x_vector_reg_5_6_inst : DFF_X1 port map( D => n239, CK => clk, Q => 
                           x_vector_56_port, QN => n315);
   x_vector_reg_6_6_inst : DFF_X1 port map( D => n238, CK => clk, Q => 
                           x_vector_66_port, QN => n365);
   x_vector_reg_7_6_inst : DFF_X1 port map( D => n237, CK => clk, Q => 
                           x_vector_76_port, QN => n314);
   x_vector_reg_8_6_inst : DFF_X1 port map( D => n236, CK => clk, Q => 
                           x_vector_86_port, QN => n372);
   x_vector_reg_9_6_inst : DFF_X1 port map( D => n235, CK => clk, Q => 
                           x_vector_96_port, QN => n308);
   x_vector_reg_10_6_inst : DFF_X1 port map( D => n234, CK => clk, Q => 
                           x_vector_106_port, QN => n394);
   x_vector_reg_0_5_inst : DFF_X1 port map( D => n233, CK => clk, Q => 
                           x_vector_5_port, QN => n358);
   x_vector_reg_1_5_inst : DFF_X1 port map( D => n232, CK => clk, Q => 
                           x_vector_15_port, QN => n301);
   x_vector_reg_2_5_inst : DFF_X1 port map( D => n231, CK => clk, Q => 
                           x_vector_25_port, QN => n353);
   x_vector_reg_3_5_inst : DFF_X1 port map( D => n230, CK => clk, Q => 
                           x_vector_35_port, QN => n300);
   x_vector_reg_4_5_inst : DFF_X1 port map( D => n229, CK => clk, Q => 
                           x_vector_45_port, QN => n352);
   x_vector_reg_5_5_inst : DFF_X1 port map( D => n228, CK => clk, Q => 
                           x_vector_55_port, QN => n299);
   x_vector_reg_6_5_inst : DFF_X1 port map( D => n227, CK => clk, Q => 
                           x_vector_65_port, QN => n351);
   x_vector_reg_7_5_inst : DFF_X1 port map( D => n226, CK => clk, Q => 
                           x_vector_75_port, QN => n298);
   x_vector_reg_8_5_inst : DFF_X1 port map( D => n225, CK => clk, Q => 
                           x_vector_85_port, QN => n350);
   x_vector_reg_9_5_inst : DFF_X1 port map( D => n224, CK => clk, Q => 
                           x_vector_95_port, QN => n306);
   x_vector_reg_10_5_inst : DFF_X1 port map( D => n223, CK => clk, Q => 
                           x_vector_105_port, QN => n390);
   x_vector_reg_0_4_inst : DFF_X1 port map( D => n222, CK => clk, Q => 
                           x_vector_4_port, QN => n377);
   x_vector_reg_1_4_inst : DFF_X1 port map( D => n221, CK => clk, Q => 
                           x_vector_14_port, QN => n320);
   x_vector_reg_2_4_inst : DFF_X1 port map( D => n220, CK => clk, Q => 
                           x_vector_24_port, QN => n371);
   x_vector_reg_3_4_inst : DFF_X1 port map( D => n219, CK => clk, Q => 
                           x_vector_34_port, QN => n319);
   x_vector_reg_4_4_inst : DFF_X1 port map( D => n218, CK => clk, Q => 
                           x_vector_44_port, QN => n370);
   x_vector_reg_5_4_inst : DFF_X1 port map( D => n217, CK => clk, Q => 
                           x_vector_54_port, QN => n318);
   x_vector_reg_6_4_inst : DFF_X1 port map( D => n216, CK => clk, Q => 
                           x_vector_64_port, QN => n369);
   x_vector_reg_7_4_inst : DFF_X1 port map( D => n215, CK => clk, Q => 
                           x_vector_74_port, QN => n317);
   x_vector_reg_8_4_inst : DFF_X1 port map( D => n214, CK => clk, Q => 
                           x_vector_84_port, QN => n368);
   x_vector_reg_9_4_inst : DFF_X1 port map( D => n213, CK => clk, Q => 
                           x_vector_94_port, QN => n326);
   x_vector_reg_10_4_inst : DFF_X1 port map( D => n212_port, CK => clk, Q => 
                           x_vector_104_port, QN => n393);
   x_vector_reg_0_3_inst : DFF_X1 port map( D => n211_port, CK => clk, Q => 
                           x_vector_3_port, QN => n348);
   x_vector_reg_1_3_inst : DFF_X1 port map( D => n210_port, CK => clk, Q => 
                           x_vector_13_port, QN => n296);
   x_vector_reg_2_3_inst : DFF_X1 port map( D => n209_port, CK => clk, Q => 
                           x_vector_23_port, QN => n347);
   x_vector_reg_3_3_inst : DFF_X1 port map( D => n208_port, CK => clk, Q => 
                           x_vector_33_port, QN => n295);
   x_vector_reg_4_3_inst : DFF_X1 port map( D => n207_port, CK => clk, Q => 
                           x_vector_43_port, QN => n346);
   x_vector_reg_5_3_inst : DFF_X1 port map( D => n206_port, CK => clk, Q => 
                           x_vector_53_port, QN => n294);
   x_vector_reg_6_3_inst : DFF_X1 port map( D => n205_port, CK => clk, Q => 
                           x_vector_63_port, QN => n345);
   x_vector_reg_7_3_inst : DFF_X1 port map( D => n204_port, CK => clk, Q => 
                           x_vector_73_port, QN => n293);
   x_vector_reg_8_3_inst : DFF_X1 port map( D => n203_port, CK => clk, Q => 
                           x_vector_83_port, QN => n344);
   x_vector_reg_9_3_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           x_vector_93_port, QN => n297);
   x_vector_reg_10_3_inst : DFF_X1 port map( D => n201, CK => clk, Q => 
                           x_vector_103_port, QN => n349);
   x_vector_reg_0_2_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           x_vector_2_port, QN => n384);
   x_vector_reg_1_2_inst : DFF_X1 port map( D => n199, CK => clk, Q => 
                           x_vector_12_port, QN => n331);
   x_vector_reg_2_2_inst : DFF_X1 port map( D => n198, CK => clk, Q => 
                           x_vector_22_port, QN => n383);
   x_vector_reg_3_2_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           x_vector_32_port, QN => n330);
   x_vector_reg_4_2_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           x_vector_42_port, QN => n382);
   x_vector_reg_5_2_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           x_vector_52_port, QN => n329);
   x_vector_reg_6_2_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           x_vector_62_port, QN => n381);
   x_vector_reg_7_2_inst : DFF_X1 port map( D => n193, CK => clk, Q => 
                           x_vector_72_port, QN => n328);
   x_vector_reg_8_2_inst : DFF_X1 port map( D => n192, CK => clk, Q => 
                           x_vector_82_port, QN => n380);
   x_vector_reg_9_2_inst : DFF_X1 port map( D => n191, CK => clk, Q => 
                           x_vector_92_port, QN => n332);
   x_vector_reg_10_2_inst : DFF_X1 port map( D => n190, CK => clk, Q => 
                           x_vector_102_port, QN => n396);
   x_vector_reg_0_1_inst : DFF_X1 port map( D => n189, CK => clk, Q => 
                           x_vector_1_port, QN => n342);
   x_vector_reg_1_1_inst : DFF_X1 port map( D => n188, CK => clk, Q => 
                           x_vector_11_port, QN => n291);
   x_vector_reg_2_1_inst : DFF_X1 port map( D => n187, CK => clk, Q => 
                           x_vector_21_port, QN => n341);
   x_vector_reg_3_1_inst : DFF_X1 port map( D => n186, CK => clk, Q => 
                           x_vector_31_port, QN => n290);
   x_vector_reg_4_1_inst : DFF_X1 port map( D => n185, CK => clk, Q => 
                           x_vector_41_port, QN => n340);
   x_vector_reg_5_1_inst : DFF_X1 port map( D => n184, CK => clk, Q => 
                           x_vector_51_port, QN => n289);
   x_vector_reg_6_1_inst : DFF_X1 port map( D => n183, CK => clk, Q => 
                           x_vector_61_port, QN => n339);
   x_vector_reg_7_1_inst : DFF_X1 port map( D => n182, CK => clk, Q => 
                           x_vector_71_port, QN => n288);
   x_vector_reg_8_1_inst : DFF_X1 port map( D => n181, CK => clk, Q => 
                           x_vector_81_port, QN => n338);
   x_vector_reg_9_1_inst : DFF_X1 port map( D => n180, CK => clk, Q => 
                           x_vector_91_port, QN => n292);
   x_vector_reg_10_1_inst : DFF_X1 port map( D => n179, CK => clk, Q => 
                           x_vector_101_port, QN => n343);
   x_vector_reg_0_0_inst : DFF_X1 port map( D => n178, CK => clk, Q => 
                           x_vector_0_port, QN => n389);
   x_vector_reg_1_0_inst : DFF_X1 port map( D => n177, CK => clk, Q => 
                           x_vector_10_port, QN => n336);
   x_vector_reg_2_0_inst : DFF_X1 port map( D => n176, CK => clk, Q => 
                           x_vector_20_port, QN => n388);
   x_vector_reg_3_0_inst : DFF_X1 port map( D => n175, CK => clk, Q => 
                           x_vector_30_port, QN => n335);
   x_vector_reg_4_0_inst : DFF_X1 port map( D => n174, CK => clk, Q => 
                           x_vector_40_port, QN => n387);
   x_vector_reg_5_0_inst : DFF_X1 port map( D => n173, CK => clk, Q => 
                           x_vector_50_port, QN => n334);
   x_vector_reg_6_0_inst : DFF_X1 port map( D => n172, CK => clk, Q => 
                           x_vector_60_port, QN => n386);
   x_vector_reg_7_0_inst : DFF_X1 port map( D => n171, CK => clk, Q => 
                           x_vector_70_port, QN => n333);
   x_vector_reg_8_0_inst : DFF_X1 port map( D => n170, CK => clk, Q => 
                           x_vector_80_port, QN => n385);
   x_vector_reg_9_0_inst : DFF_X1 port map( D => n169, CK => clk, Q => 
                           x_vector_90_port, QN => n337);
   x_vector_reg_10_0_inst : DFF_X1 port map( D => n168, CK => clk, Q => 
                           x_vector_100_port, QN => n397);
   VOUT_reg : DFF_X1 port map( D => n167, CK => clk, Q => VOUT, QN => n156);
   U259 : BUF_X1 port map( A => n410, Z => n413);
   U260 : BUF_X1 port map( A => n411, Z => n416);
   U261 : BUF_X1 port map( A => n411, Z => n417);
   U262 : BUF_X1 port map( A => n410, Z => n415);
   U263 : BUF_X1 port map( A => n410, Z => n414);
   U264 : BUF_X1 port map( A => n411, Z => n418);
   U265 : BUF_X1 port map( A => n412, Z => n420);
   U266 : BUF_X1 port map( A => n412, Z => n419);
   U267 : BUF_X1 port map( A => n398, Z => n404);
   U268 : BUF_X1 port map( A => n398, Z => n405);
   U269 : BUF_X1 port map( A => n398, Z => n400);
   U270 : BUF_X1 port map( A => n398, Z => n401);
   U271 : BUF_X1 port map( A => n398, Z => n402);
   U272 : BUF_X1 port map( A => n398, Z => n403);
   U273 : BUF_X1 port map( A => n399, Z => n406);
   U274 : BUF_X1 port map( A => n399, Z => n407);
   U275 : BUF_X1 port map( A => n399, Z => n408);
   U276 : OAI22_X1 port map( A1 => n421, A2 => n372, B1 => n400, B2 => n314, ZN
                           => n236);
   U277 : OAI22_X1 port map( A1 => n421, A2 => n314, B1 => n400, B2 => n365, ZN
                           => n237);
   U278 : OAI22_X1 port map( A1 => n421, A2 => n365, B1 => n400, B2 => n315, ZN
                           => n238);
   U279 : OAI22_X1 port map( A1 => n421, A2 => n315, B1 => n400, B2 => n366, ZN
                           => n239);
   U280 : OAI22_X1 port map( A1 => n421, A2 => n366, B1 => n400, B2 => n316, ZN
                           => n240);
   U281 : OAI22_X1 port map( A1 => n421, A2 => n316, B1 => n400, B2 => n367, ZN
                           => n241);
   U282 : OAI22_X1 port map( A1 => n421, A2 => n367, B1 => n400, B2 => n321, ZN
                           => n242);
   U283 : OAI22_X1 port map( A1 => n417, A2 => n292, B1 => n404, B2 => n338, ZN
                           => n180);
   U284 : OAI22_X1 port map( A1 => n417, A2 => n338, B1 => n404, B2 => n288, ZN
                           => n181);
   U285 : OAI22_X1 port map( A1 => n417, A2 => n288, B1 => n404, B2 => n339, ZN
                           => n182);
   U286 : OAI22_X1 port map( A1 => n417, A2 => n339, B1 => n404, B2 => n289, ZN
                           => n183);
   U287 : OAI22_X1 port map( A1 => n416, A2 => n289, B1 => n405, B2 => n340, ZN
                           => n184);
   U288 : OAI22_X1 port map( A1 => n416, A2 => n340, B1 => n405, B2 => n290, ZN
                           => n185);
   U289 : OAI22_X1 port map( A1 => n416, A2 => n290, B1 => n405, B2 => n341, ZN
                           => n186);
   U290 : OAI22_X1 port map( A1 => n416, A2 => n341, B1 => n405, B2 => n291, ZN
                           => n187);
   U291 : OAI22_X1 port map( A1 => n416, A2 => n291, B1 => n405, B2 => n342, ZN
                           => n188);
   U292 : OAI22_X1 port map( A1 => n415, A2 => n297, B1 => n406, B2 => n344, ZN
                           => n202);
   U293 : OAI22_X1 port map( A1 => n415, A2 => n344, B1 => n406, B2 => n293, ZN
                           => n203_port);
   U294 : OAI22_X1 port map( A1 => n415, A2 => n293, B1 => n406, B2 => n345, ZN
                           => n204_port);
   U295 : OAI22_X1 port map( A1 => n415, A2 => n345, B1 => n406, B2 => n294, ZN
                           => n205_port);
   U296 : OAI22_X1 port map( A1 => n415, A2 => n294, B1 => n406, B2 => n346, ZN
                           => n206_port);
   U297 : OAI22_X1 port map( A1 => n415, A2 => n346, B1 => n406, B2 => n295, ZN
                           => n207_port);
   U298 : OAI22_X1 port map( A1 => n417, A2 => n295, B1 => n407, B2 => n347, ZN
                           => n208_port);
   U299 : OAI22_X1 port map( A1 => n415, A2 => n347, B1 => n407, B2 => n296, ZN
                           => n209_port);
   U300 : OAI22_X1 port map( A1 => n415, A2 => n296, B1 => n407, B2 => n348, ZN
                           => n210_port);
   U301 : OAI22_X1 port map( A1 => n418, A2 => n337, B1 => n403, B2 => n385, ZN
                           => n169);
   U302 : OAI22_X1 port map( A1 => n418, A2 => n385, B1 => n403, B2 => n333, ZN
                           => n170);
   U303 : OAI22_X1 port map( A1 => n418, A2 => n333, B1 => n403, B2 => n386, ZN
                           => n171);
   U304 : OAI22_X1 port map( A1 => n417, A2 => n386, B1 => n404, B2 => n334, ZN
                           => n172);
   U305 : OAI22_X1 port map( A1 => n417, A2 => n334, B1 => n404, B2 => n387, ZN
                           => n173);
   U306 : OAI22_X1 port map( A1 => n417, A2 => n387, B1 => n404, B2 => n335, ZN
                           => n174);
   U307 : OAI22_X1 port map( A1 => n417, A2 => n335, B1 => n404, B2 => n388, ZN
                           => n175);
   U308 : OAI22_X1 port map( A1 => n417, A2 => n388, B1 => n404, B2 => n336, ZN
                           => n176);
   U309 : OAI22_X1 port map( A1 => n417, A2 => n336, B1 => n404, B2 => n389, ZN
                           => n177);
   U310 : OAI22_X1 port map( A1 => n416, A2 => n332, B1 => n405, B2 => n380, ZN
                           => n191);
   U311 : OAI22_X1 port map( A1 => n416, A2 => n380, B1 => n405, B2 => n328, ZN
                           => n192);
   U312 : OAI22_X1 port map( A1 => n416, A2 => n328, B1 => n405, B2 => n381, ZN
                           => n193);
   U313 : OAI22_X1 port map( A1 => n416, A2 => n381, B1 => n405, B2 => n329, ZN
                           => n194);
   U314 : OAI22_X1 port map( A1 => n416, A2 => n329, B1 => n405, B2 => n382, ZN
                           => n195);
   U315 : OAI22_X1 port map( A1 => n416, A2 => n382, B1 => n406, B2 => n330, ZN
                           => n196);
   U316 : OAI22_X1 port map( A1 => n415, A2 => n330, B1 => n406, B2 => n383, ZN
                           => n197);
   U317 : OAI22_X1 port map( A1 => n415, A2 => n383, B1 => n406, B2 => n331, ZN
                           => n198);
   U318 : OAI22_X1 port map( A1 => n415, A2 => n331, B1 => n406, B2 => n384, ZN
                           => n199);
   U319 : OAI22_X1 port map( A1 => n414, A2 => n326, B1 => n407, B2 => n368, ZN
                           => n213);
   U320 : OAI22_X1 port map( A1 => n414, A2 => n368, B1 => n407, B2 => n317, ZN
                           => n214);
   U321 : OAI22_X1 port map( A1 => n414, A2 => n317, B1 => n407, B2 => n369, ZN
                           => n215);
   U322 : OAI22_X1 port map( A1 => n414, A2 => n369, B1 => n407, B2 => n318, ZN
                           => n216);
   U323 : OAI22_X1 port map( A1 => n414, A2 => n318, B1 => n407, B2 => n370, ZN
                           => n217);
   U324 : OAI22_X1 port map( A1 => n414, A2 => n370, B1 => n407, B2 => n319, ZN
                           => n218);
   U325 : OAI22_X1 port map( A1 => n414, A2 => n319, B1 => n407, B2 => n371, ZN
                           => n219);
   U326 : OAI22_X1 port map( A1 => n414, A2 => n371, B1 => n408, B2 => n320, ZN
                           => n220);
   U327 : OAI22_X1 port map( A1 => n414, A2 => n320, B1 => n408, B2 => n377, ZN
                           => n221);
   U328 : OAI22_X1 port map( A1 => n308, A2 => n413, B1 => n400, B2 => n372, ZN
                           => n235);
   U329 : OAI22_X1 port map( A1 => n420, A2 => n321, B1 => n400, B2 => n378, ZN
                           => n243);
   U330 : OAI22_X1 port map( A1 => n419, A2 => n327, B1 => n401, B2 => n373, ZN
                           => n257);
   U331 : OAI22_X1 port map( A1 => n419, A2 => n373, B1 => n402, B2 => n322, ZN
                           => n258);
   U332 : OAI22_X1 port map( A1 => n419, A2 => n322, B1 => n402, B2 => n374, ZN
                           => n259);
   U333 : OAI22_X1 port map( A1 => n419, A2 => n374, B1 => n402, B2 => n323, ZN
                           => n260);
   U334 : OAI22_X1 port map( A1 => n419, A2 => n323, B1 => n402, B2 => n375, ZN
                           => n261);
   U335 : OAI22_X1 port map( A1 => n419, A2 => n375, B1 => n402, B2 => n324, ZN
                           => n262);
   U336 : OAI22_X1 port map( A1 => n419, A2 => n324, B1 => n402, B2 => n376, ZN
                           => n263);
   U337 : OAI22_X1 port map( A1 => n419, A2 => n376, B1 => n402, B2 => n325, ZN
                           => n264);
   U338 : OAI22_X1 port map( A1 => n419, A2 => n325, B1 => n402, B2 => n379, ZN
                           => n265);
   U339 : OAI22_X1 port map( A1 => n419, A2 => n313, B1 => n402, B2 => n360, ZN
                           => n268);
   U340 : OAI22_X1 port map( A1 => n418, A2 => n360, B1 => n402, B2 => n309, ZN
                           => n269);
   U341 : OAI22_X1 port map( A1 => n418, A2 => n309, B1 => n403, B2 => n361, ZN
                           => n270);
   U342 : OAI22_X1 port map( A1 => n418, A2 => n361, B1 => n403, B2 => n310, ZN
                           => n271);
   U343 : OAI22_X1 port map( A1 => n418, A2 => n310, B1 => n403, B2 => n362, ZN
                           => n272);
   U344 : OAI22_X1 port map( A1 => n418, A2 => n362, B1 => n403, B2 => n311, ZN
                           => n273);
   U345 : OAI22_X1 port map( A1 => n418, A2 => n311, B1 => n403, B2 => n363, ZN
                           => n274);
   U346 : OAI22_X1 port map( A1 => n418, A2 => n363, B1 => n403, B2 => n312, ZN
                           => n275);
   U347 : OAI22_X1 port map( A1 => n418, A2 => n312, B1 => n403, B2 => n364, ZN
                           => n276);
   U348 : OAI22_X1 port map( A1 => n414, A2 => n306, B1 => n408, B2 => n350, ZN
                           => n224);
   U349 : OAI22_X1 port map( A1 => n413, A2 => n350, B1 => n408, B2 => n298, ZN
                           => n225);
   U350 : OAI22_X1 port map( A1 => n413, A2 => n298, B1 => n408, B2 => n351, ZN
                           => n226);
   U351 : OAI22_X1 port map( A1 => n413, A2 => n351, B1 => n408, B2 => n299, ZN
                           => n227);
   U352 : OAI22_X1 port map( A1 => n413, A2 => n299, B1 => n408, B2 => n352, ZN
                           => n228);
   U353 : OAI22_X1 port map( A1 => n413, A2 => n352, B1 => n408, B2 => n300, ZN
                           => n229);
   U354 : OAI22_X1 port map( A1 => n413, A2 => n300, B1 => n408, B2 => n353, ZN
                           => n230);
   U355 : OAI22_X1 port map( A1 => n413, A2 => n353, B1 => n408, B2 => n301, ZN
                           => n231);
   U356 : OAI22_X1 port map( A1 => n413, A2 => n301, B1 => n409, B2 => n358, ZN
                           => n232);
   U357 : OAI22_X1 port map( A1 => n420, A2 => n307, B1 => n401, B2 => n354, ZN
                           => n246);
   U358 : OAI22_X1 port map( A1 => n420, A2 => n354, B1 => n401, B2 => n302, ZN
                           => n247);
   U359 : OAI22_X1 port map( A1 => n420, A2 => n302, B1 => n401, B2 => n355, ZN
                           => n248);
   U360 : OAI22_X1 port map( A1 => n420, A2 => n355, B1 => n401, B2 => n303, ZN
                           => n249);
   U361 : OAI22_X1 port map( A1 => n420, A2 => n303, B1 => n401, B2 => n356, ZN
                           => n250);
   U362 : OAI22_X1 port map( A1 => n420, A2 => n356, B1 => n401, B2 => n304, ZN
                           => n251);
   U363 : OAI22_X1 port map( A1 => n420, A2 => n304, B1 => n401, B2 => n357, ZN
                           => n252);
   U364 : OAI22_X1 port map( A1 => n420, A2 => n357, B1 => n401, B2 => n305, ZN
                           => n253);
   U365 : OAI22_X1 port map( A1 => n420, A2 => n305, B1 => n401, B2 => n359, ZN
                           => n254);
   U366 : INV_X1 port map( A => n72, ZN => n443);
   U367 : BUF_X1 port map( A => n23, Z => n398);
   U368 : BUF_X1 port map( A => n23, Z => n399);
   U369 : OAI22_X1 port map( A1 => n158, A2 => n443, B1 => n72, B2 => n430, ZN 
                           => n279);
   U370 : INV_X1 port map( A => N204, ZN => n430);
   U371 : OAI22_X1 port map( A1 => n159, A2 => n443, B1 => n72, B2 => n429, ZN 
                           => n280);
   U372 : INV_X1 port map( A => N205, ZN => n429);
   U373 : OAI22_X1 port map( A1 => n161, A2 => n443, B1 => n72, B2 => n427, ZN 
                           => n282);
   U374 : INV_X1 port map( A => N207, ZN => n427);
   U375 : OAI22_X1 port map( A1 => n162, A2 => n443, B1 => n72, B2 => n426, ZN 
                           => n283);
   U376 : INV_X1 port map( A => N208, ZN => n426);
   U377 : OAI22_X1 port map( A1 => n163, A2 => n443, B1 => n72, B2 => n425, ZN 
                           => n284);
   U378 : INV_X1 port map( A => N209, ZN => n425);
   U379 : OAI22_X1 port map( A1 => n164, A2 => n443, B1 => n72, B2 => n424, ZN 
                           => n285);
   U380 : INV_X1 port map( A => N210, ZN => n424);
   U381 : OAI22_X1 port map( A1 => n165, A2 => n443, B1 => n72, B2 => n423, ZN 
                           => n286);
   U382 : INV_X1 port map( A => N211, ZN => n423);
   U383 : OAI22_X1 port map( A1 => n160, A2 => n443, B1 => n72, B2 => n428, ZN 
                           => n281);
   U384 : INV_X1 port map( A => N206, ZN => n428);
   U385 : OAI22_X1 port map( A1 => n166, A2 => n443, B1 => n72, B2 => n422, ZN 
                           => n287);
   U386 : INV_X1 port map( A => N212, ZN => n422);
   U387 : OAI22_X1 port map( A1 => n157, A2 => n443, B1 => n72, B2 => n431, ZN 
                           => n278);
   U388 : INV_X1 port map( A => N203, ZN => n431);
   U389 : OAI22_X1 port map( A1 => n417, A2 => n343, B1 => n404, B2 => n292, ZN
                           => n179);
   U390 : OAI22_X1 port map( A1 => n415, A2 => n349, B1 => n406, B2 => n297, ZN
                           => n201);
   U391 : OAI22_X1 port map( A1 => n417, A2 => n389, B1 => n404, B2 => n441, ZN
                           => n178);
   U392 : INV_X1 port map( A => DIN(0), ZN => n441);
   U393 : OAI22_X1 port map( A1 => n416, A2 => n342, B1 => n405, B2 => n440, ZN
                           => n189);
   U394 : INV_X1 port map( A => DIN(1), ZN => n440);
   U395 : OAI22_X1 port map( A1 => n415, A2 => n384, B1 => n406, B2 => n439, ZN
                           => n200);
   U396 : INV_X1 port map( A => DIN(2), ZN => n439);
   U397 : OAI22_X1 port map( A1 => n414, A2 => n348, B1 => n407, B2 => n438, ZN
                           => n211_port);
   U398 : INV_X1 port map( A => DIN(3), ZN => n438);
   U399 : OAI22_X1 port map( A1 => n414, A2 => n377, B1 => n408, B2 => n437, ZN
                           => n222);
   U400 : INV_X1 port map( A => DIN(4), ZN => n437);
   U401 : OAI22_X1 port map( A1 => n413, A2 => n358, B1 => n409, B2 => n436, ZN
                           => n233);
   U402 : INV_X1 port map( A => DIN(5), ZN => n436);
   U403 : OAI22_X1 port map( A1 => n420, A2 => n378, B1 => n400, B2 => n435, ZN
                           => n244);
   U404 : INV_X1 port map( A => DIN(6), ZN => n435);
   U405 : OAI22_X1 port map( A1 => n420, A2 => n359, B1 => n401, B2 => n434, ZN
                           => n255);
   U406 : INV_X1 port map( A => DIN(7), ZN => n434);
   U407 : OAI22_X1 port map( A1 => n419, A2 => n379, B1 => n402, B2 => n433, ZN
                           => n266);
   U408 : INV_X1 port map( A => DIN(8), ZN => n433);
   U409 : OAI22_X1 port map( A1 => n418, A2 => n364, B1 => n403, B2 => n432, ZN
                           => n277);
   U410 : INV_X1 port map( A => DIN(9), ZN => n432);
   U411 : OAI22_X1 port map( A1 => n418, A2 => n397, B1 => n403, B2 => n337, ZN
                           => n168);
   U412 : OAI22_X1 port map( A1 => n416, A2 => n396, B1 => n405, B2 => n332, ZN
                           => n190);
   U413 : OAI22_X1 port map( A1 => n414, A2 => n393, B1 => n407, B2 => n326, ZN
                           => n212_port);
   U414 : OAI22_X1 port map( A1 => n413, A2 => n394, B1 => n400, B2 => n308, ZN
                           => n234);
   U415 : OAI22_X1 port map( A1 => n419, A2 => n395, B1 => n401, B2 => n327, ZN
                           => n256);
   U416 : OAI22_X1 port map( A1 => n419, A2 => n392, B1 => n402, B2 => n313, ZN
                           => n267);
   U417 : OAI22_X1 port map( A1 => n413, A2 => n390, B1 => n408, B2 => n306, ZN
                           => n223);
   U418 : OAI22_X1 port map( A1 => n420, A2 => n391, B1 => n400, B2 => n307, ZN
                           => n245);
   U419 : OAI21_X1 port map( B1 => rst_n, B2 => n156, A => n72, ZN => n167);
   U420 : NAND2_X1 port map( A1 => VIN, A2 => rst_n, ZN => n72);
   U421 : NAND2_X1 port map( A1 => rst_n, A2 => n413, ZN => n23);
   U422 : NAND2_X1 port map( A1 => rst_n, A2 => n442, ZN => n21);
   U423 : INV_X1 port map( A => VIN, ZN => n442);
   U424 : CLKBUF_X1 port map( A => n399, Z => n409);
   U425 : CLKBUF_X1 port map( A => n21, Z => n410);
   U426 : CLKBUF_X1 port map( A => n21, Z => n411);
   U427 : CLKBUF_X1 port map( A => n21, Z => n412);
   U428 : CLKBUF_X1 port map( A => n412, Z => n421);
   n444 <= '0';
   n445 <= '0';
   n446 <= '0';
   n447 <= '0';
   n448 <= '0';
   n449 <= '0';
   n450 <= '0';
   n451 <= '0';
   n452 <= '0';
   n453 <= '0';
   mult_42_U391 : NAND2_X1 port map( A1 => x_vector_1_port, A2 => mult_42_n320,
                           ZN => mult_42_n341);
   mult_42_U390 : XNOR2_X1 port map( A => B(2), B => x_vector_1_port, ZN => 
                           mult_42_n340);
   mult_42_U389 : OAI22_X1 port map( A1 => B(1), A2 => mult_42_n341, B1 => 
                           mult_42_n340, B2 => mult_42_n320, ZN => mult_42_n402
                           );
   mult_42_U388 : NAND3_X1 port map( A1 => mult_42_n402, A2 => mult_42_n312, A3
                           => x_vector_1_port, ZN => mult_42_n400);
   mult_42_U387 : XNOR2_X1 port map( A => x_vector_2_port, B => x_vector_1_port
                           , ZN => mult_42_n352);
   mult_42_U386 : NAND2_X1 port map( A1 => mult_42_n319, A2 => mult_42_n402, ZN
                           => mult_42_n401);
   mult_42_U385 : MUX2_X1 port map( A => mult_42_n400, B => mult_42_n401, S => 
                           B(0), Z => mult_42_n396);
   mult_42_U384 : XOR2_X1 port map( A => x_vector_3_port, B => x_vector_2_port,
                           Z => mult_42_n399);
   mult_42_U383 : NAND2_X1 port map( A1 => mult_42_n352, A2 => mult_42_n399, ZN
                           => mult_42_n351);
   mult_42_U382 : NOR3_X1 port map( A1 => mult_42_n352, A2 => B(0), A3 => 
                           mult_42_n317, ZN => mult_42_n398);
   mult_42_U381 : AOI21_X1 port map( B1 => x_vector_3_port, B2 => mult_42_n318,
                           A => mult_42_n398, ZN => mult_42_n397);
   mult_42_U380 : OAI222_X1 port map( A1 => mult_42_n396, A2 => mult_42_n311, 
                           B1 => mult_42_n397, B2 => mult_42_n396, C1 => 
                           mult_42_n397, C2 => mult_42_n311, ZN => mult_42_n395
                           );
   mult_42_U379 : AOI222_X1 port map( A1 => mult_42_n395, A2 => mult_42_n88, B1
                           => mult_42_n395, B2 => mult_42_n89, C1 => 
                           mult_42_n89, C2 => mult_42_n88, ZN => mult_42_n394);
   mult_42_U378 : OAI222_X1 port map( A1 => mult_42_n394, A2 => mult_42_n308, 
                           B1 => mult_42_n394, B2 => mult_42_n309, C1 => 
                           mult_42_n309, C2 => mult_42_n308, ZN => mult_42_n393
                           );
   mult_42_U377 : AOI222_X1 port map( A1 => mult_42_n393, A2 => mult_42_n80, B1
                           => mult_42_n393, B2 => mult_42_n83, C1 => 
                           mult_42_n83, C2 => mult_42_n80, ZN => mult_42_n392);
   mult_42_U376 : OAI222_X1 port map( A1 => mult_42_n392, A2 => mult_42_n305, 
                           B1 => mult_42_n392, B2 => mult_42_n307, C1 => 
                           mult_42_n307, C2 => mult_42_n305, ZN => mult_42_n391
                           );
   mult_42_U375 : AOI222_X1 port map( A1 => mult_42_n391, A2 => mult_42_n68, B1
                           => mult_42_n391, B2 => mult_42_n73, C1 => 
                           mult_42_n73, C2 => mult_42_n68, ZN => mult_42_n390);
   mult_42_U374 : OAI222_X1 port map( A1 => mult_42_n390, A2 => mult_42_n296, 
                           B1 => mult_42_n390, B2 => mult_42_n304, C1 => 
                           mult_42_n304, C2 => mult_42_n296, ZN => mult_42_n10)
                           ;
   mult_42_U373 : XOR2_X1 port map( A => x_vector_9_port, B => x_vector_8_port,
                           Z => mult_42_n389);
   mult_42_U372 : NAND2_X1 port map( A1 => mult_42_n338, A2 => mult_42_n389, ZN
                           => mult_42_n337);
   mult_42_U371 : OR3_X1 port map( A1 => mult_42_n338, A2 => B(0), A3 => 
                           mult_42_n314, ZN => mult_42_n388);
   mult_42_U370 : OAI21_X1 port map( B1 => mult_42_n314, B2 => mult_42_n337, A 
                           => mult_42_n388, ZN => mult_42_n105);
   mult_42_U369 : XOR2_X1 port map( A => x_vector_7_port, B => x_vector_6_port,
                           Z => mult_42_n387);
   mult_42_U368 : NAND2_X1 port map( A1 => mult_42_n327, A2 => mult_42_n387, ZN
                           => mult_42_n326);
   mult_42_U367 : OR3_X1 port map( A1 => mult_42_n327, A2 => B(0), A3 => 
                           mult_42_n315, ZN => mult_42_n386);
   mult_42_U366 : OAI21_X1 port map( B1 => mult_42_n315, B2 => mult_42_n326, A 
                           => mult_42_n386, ZN => mult_42_n106);
   mult_42_U365 : XOR2_X1 port map( A => x_vector_5_port, B => x_vector_4_port,
                           Z => mult_42_n385);
   mult_42_U364 : NAND2_X1 port map( A1 => mult_42_n332, A2 => mult_42_n385, ZN
                           => mult_42_n331);
   mult_42_U363 : OR3_X1 port map( A1 => mult_42_n332, A2 => B(0), A3 => 
                           mult_42_n316, ZN => mult_42_n384);
   mult_42_U362 : OAI21_X1 port map( B1 => mult_42_n316, B2 => mult_42_n331, A 
                           => mult_42_n384, ZN => mult_42_n107);
   mult_42_U361 : XOR2_X1 port map( A => B(9), B => mult_42_n314, Z => 
                           mult_42_n339);
   mult_42_U360 : OAI22_X1 port map( A1 => mult_42_n339, A2 => mult_42_n338, B1
                           => mult_42_n337, B2 => mult_42_n339, ZN => 
                           mult_42_n383);
   mult_42_U359 : XOR2_X1 port map( A => B(7), B => mult_42_n314, Z => 
                           mult_42_n382);
   mult_42_U358 : XOR2_X1 port map( A => B(8), B => mult_42_n314, Z => 
                           mult_42_n336);
   mult_42_U357 : OAI22_X1 port map( A1 => mult_42_n382, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n336, ZN => 
                           mult_42_n111);
   mult_42_U356 : XOR2_X1 port map( A => B(6), B => mult_42_n314, Z => 
                           mult_42_n381);
   mult_42_U355 : OAI22_X1 port map( A1 => mult_42_n381, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n382, ZN => 
                           mult_42_n112);
   mult_42_U354 : XOR2_X1 port map( A => B(5), B => mult_42_n314, Z => 
                           mult_42_n380);
   mult_42_U353 : OAI22_X1 port map( A1 => mult_42_n380, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n381, ZN => 
                           mult_42_n113);
   mult_42_U352 : XOR2_X1 port map( A => B(4), B => mult_42_n314, Z => 
                           mult_42_n379);
   mult_42_U351 : OAI22_X1 port map( A1 => mult_42_n379, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n380, ZN => 
                           mult_42_n114);
   mult_42_U350 : XOR2_X1 port map( A => B(3), B => mult_42_n314, Z => 
                           mult_42_n378);
   mult_42_U349 : OAI22_X1 port map( A1 => mult_42_n378, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n379, ZN => 
                           mult_42_n115);
   mult_42_U348 : XOR2_X1 port map( A => B(2), B => mult_42_n314, Z => 
                           mult_42_n377);
   mult_42_U347 : OAI22_X1 port map( A1 => mult_42_n377, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n378, ZN => 
                           mult_42_n116);
   mult_42_U346 : XOR2_X1 port map( A => mult_42_n312, B => x_vector_9_port, Z 
                           => mult_42_n376);
   mult_42_U345 : OAI22_X1 port map( A1 => mult_42_n376, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n377, ZN => 
                           mult_42_n117);
   mult_42_U344 : XOR2_X1 port map( A => mult_42_n314, B => B(0), Z => 
                           mult_42_n375);
   mult_42_U343 : OAI22_X1 port map( A1 => mult_42_n375, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n376, ZN => 
                           mult_42_n118);
   mult_42_U342 : NOR2_X1 port map( A1 => mult_42_n338, A2 => mult_42_n313, ZN 
                           => mult_42_n119);
   mult_42_U341 : XOR2_X1 port map( A => B(9), B => mult_42_n315, Z => 
                           mult_42_n335);
   mult_42_U340 : OAI22_X1 port map( A1 => mult_42_n335, A2 => mult_42_n327, B1
                           => mult_42_n326, B2 => mult_42_n335, ZN => 
                           mult_42_n374);
   mult_42_U339 : XOR2_X1 port map( A => B(7), B => mult_42_n315, Z => 
                           mult_42_n373);
   mult_42_U338 : XOR2_X1 port map( A => B(8), B => mult_42_n315, Z => 
                           mult_42_n334);
   mult_42_U337 : OAI22_X1 port map( A1 => mult_42_n373, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n334, ZN => 
                           mult_42_n121);
   mult_42_U336 : XOR2_X1 port map( A => B(6), B => mult_42_n315, Z => 
                           mult_42_n372);
   mult_42_U335 : OAI22_X1 port map( A1 => mult_42_n372, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n373, ZN => 
                           mult_42_n122);
   mult_42_U334 : XOR2_X1 port map( A => B(5), B => mult_42_n315, Z => 
                           mult_42_n371);
   mult_42_U333 : OAI22_X1 port map( A1 => mult_42_n371, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n372, ZN => 
                           mult_42_n123);
   mult_42_U332 : XOR2_X1 port map( A => B(4), B => mult_42_n315, Z => 
                           mult_42_n328);
   mult_42_U331 : OAI22_X1 port map( A1 => mult_42_n328, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n371, ZN => 
                           mult_42_n124);
   mult_42_U330 : XOR2_X1 port map( A => B(2), B => mult_42_n315, Z => 
                           mult_42_n370);
   mult_42_U329 : XOR2_X1 port map( A => B(3), B => mult_42_n315, Z => 
                           mult_42_n325);
   mult_42_U328 : OAI22_X1 port map( A1 => mult_42_n370, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n325, ZN => 
                           mult_42_n126);
   mult_42_U327 : XOR2_X1 port map( A => mult_42_n312, B => x_vector_7_port, Z 
                           => mult_42_n369);
   mult_42_U326 : OAI22_X1 port map( A1 => mult_42_n369, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n370, ZN => 
                           mult_42_n127);
   mult_42_U325 : XOR2_X1 port map( A => mult_42_n313, B => x_vector_7_port, Z 
                           => mult_42_n368);
   mult_42_U324 : OAI22_X1 port map( A1 => mult_42_n368, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n369, ZN => 
                           mult_42_n128);
   mult_42_U323 : NOR2_X1 port map( A1 => mult_42_n327, A2 => mult_42_n313, ZN 
                           => mult_42_n129);
   mult_42_U322 : XOR2_X1 port map( A => B(9), B => mult_42_n316, Z => 
                           mult_42_n333);
   mult_42_U321 : OAI22_X1 port map( A1 => mult_42_n333, A2 => mult_42_n332, B1
                           => mult_42_n331, B2 => mult_42_n333, ZN => 
                           mult_42_n367);
   mult_42_U320 : XOR2_X1 port map( A => B(7), B => mult_42_n316, Z => 
                           mult_42_n366);
   mult_42_U319 : XOR2_X1 port map( A => B(8), B => mult_42_n316, Z => 
                           mult_42_n330);
   mult_42_U318 : OAI22_X1 port map( A1 => mult_42_n366, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n330, ZN => 
                           mult_42_n131);
   mult_42_U317 : XOR2_X1 port map( A => B(6), B => mult_42_n316, Z => 
                           mult_42_n365);
   mult_42_U316 : OAI22_X1 port map( A1 => mult_42_n365, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n366, ZN => 
                           mult_42_n132);
   mult_42_U315 : XOR2_X1 port map( A => B(5), B => mult_42_n316, Z => 
                           mult_42_n364);
   mult_42_U314 : OAI22_X1 port map( A1 => mult_42_n364, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n365, ZN => 
                           mult_42_n133);
   mult_42_U313 : XOR2_X1 port map( A => B(4), B => mult_42_n316, Z => 
                           mult_42_n363);
   mult_42_U312 : OAI22_X1 port map( A1 => mult_42_n363, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n364, ZN => 
                           mult_42_n134);
   mult_42_U311 : XOR2_X1 port map( A => B(3), B => mult_42_n316, Z => 
                           mult_42_n362);
   mult_42_U310 : OAI22_X1 port map( A1 => mult_42_n362, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n363, ZN => 
                           mult_42_n135);
   mult_42_U309 : XOR2_X1 port map( A => B(2), B => mult_42_n316, Z => 
                           mult_42_n361);
   mult_42_U308 : OAI22_X1 port map( A1 => mult_42_n361, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n362, ZN => 
                           mult_42_n136);
   mult_42_U307 : XOR2_X1 port map( A => mult_42_n312, B => x_vector_5_port, Z 
                           => mult_42_n360);
   mult_42_U306 : OAI22_X1 port map( A1 => mult_42_n360, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n361, ZN => 
                           mult_42_n137);
   mult_42_U305 : XOR2_X1 port map( A => mult_42_n313, B => x_vector_5_port, Z 
                           => mult_42_n359);
   mult_42_U304 : OAI22_X1 port map( A1 => mult_42_n359, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n360, ZN => 
                           mult_42_n138);
   mult_42_U303 : NOR2_X1 port map( A1 => mult_42_n332, A2 => mult_42_n313, ZN 
                           => mult_42_n139);
   mult_42_U302 : XOR2_X1 port map( A => B(9), B => x_vector_3_port, Z => 
                           mult_42_n329);
   mult_42_U301 : AOI22_X1 port map( A1 => mult_42_n329, A2 => mult_42_n319, B1
                           => mult_42_n318, B2 => mult_42_n329, ZN => 
                           mult_42_n140);
   mult_42_U300 : XOR2_X1 port map( A => B(6), B => mult_42_n317, Z => 
                           mult_42_n358);
   mult_42_U299 : XOR2_X1 port map( A => B(7), B => mult_42_n317, Z => 
                           mult_42_n324);
   mult_42_U298 : OAI22_X1 port map( A1 => mult_42_n358, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n324, ZN => 
                           mult_42_n142);
   mult_42_U297 : XOR2_X1 port map( A => B(5), B => mult_42_n317, Z => 
                           mult_42_n357);
   mult_42_U296 : OAI22_X1 port map( A1 => mult_42_n357, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n358, ZN => 
                           mult_42_n143);
   mult_42_U295 : XOR2_X1 port map( A => B(4), B => mult_42_n317, Z => 
                           mult_42_n356);
   mult_42_U294 : OAI22_X1 port map( A1 => mult_42_n356, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n357, ZN => 
                           mult_42_n144);
   mult_42_U293 : XOR2_X1 port map( A => B(3), B => mult_42_n317, Z => 
                           mult_42_n355);
   mult_42_U292 : OAI22_X1 port map( A1 => mult_42_n355, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n356, ZN => 
                           mult_42_n145);
   mult_42_U291 : XOR2_X1 port map( A => B(2), B => mult_42_n317, Z => 
                           mult_42_n354);
   mult_42_U290 : OAI22_X1 port map( A1 => mult_42_n354, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n355, ZN => 
                           mult_42_n146);
   mult_42_U289 : XOR2_X1 port map( A => mult_42_n312, B => x_vector_3_port, Z 
                           => mult_42_n353);
   mult_42_U288 : OAI22_X1 port map( A1 => mult_42_n353, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n354, ZN => 
                           mult_42_n147);
   mult_42_U287 : XOR2_X1 port map( A => mult_42_n313, B => x_vector_3_port, Z 
                           => mult_42_n350);
   mult_42_U286 : OAI22_X1 port map( A1 => mult_42_n350, A2 => mult_42_n351, B1
                           => mult_42_n352, B2 => mult_42_n353, ZN => 
                           mult_42_n148);
   mult_42_U285 : XNOR2_X1 port map( A => B(9), B => x_vector_1_port, ZN => 
                           mult_42_n348);
   mult_42_U284 : OAI22_X1 port map( A1 => mult_42_n320, A2 => mult_42_n348, B1
                           => mult_42_n341, B2 => mult_42_n348, ZN => 
                           mult_42_n349);
   mult_42_U283 : XNOR2_X1 port map( A => B(8), B => x_vector_1_port, ZN => 
                           mult_42_n347);
   mult_42_U282 : OAI22_X1 port map( A1 => mult_42_n347, A2 => mult_42_n341, B1
                           => mult_42_n348, B2 => mult_42_n320, ZN => 
                           mult_42_n151);
   mult_42_U281 : XNOR2_X1 port map( A => B(7), B => x_vector_1_port, ZN => 
                           mult_42_n346);
   mult_42_U280 : OAI22_X1 port map( A1 => mult_42_n346, A2 => mult_42_n341, B1
                           => mult_42_n347, B2 => mult_42_n320, ZN => 
                           mult_42_n152);
   mult_42_U279 : XNOR2_X1 port map( A => B(6), B => x_vector_1_port, ZN => 
                           mult_42_n345);
   mult_42_U278 : OAI22_X1 port map( A1 => mult_42_n345, A2 => mult_42_n341, B1
                           => mult_42_n346, B2 => mult_42_n320, ZN => 
                           mult_42_n153);
   mult_42_U277 : XNOR2_X1 port map( A => B(5), B => x_vector_1_port, ZN => 
                           mult_42_n344);
   mult_42_U276 : OAI22_X1 port map( A1 => mult_42_n344, A2 => mult_42_n341, B1
                           => mult_42_n345, B2 => mult_42_n320, ZN => 
                           mult_42_n154);
   mult_42_U275 : XNOR2_X1 port map( A => B(4), B => x_vector_1_port, ZN => 
                           mult_42_n343);
   mult_42_U274 : OAI22_X1 port map( A1 => mult_42_n343, A2 => mult_42_n341, B1
                           => mult_42_n344, B2 => mult_42_n320, ZN => 
                           mult_42_n155);
   mult_42_U273 : XNOR2_X1 port map( A => B(3), B => x_vector_1_port, ZN => 
                           mult_42_n342);
   mult_42_U272 : OAI22_X1 port map( A1 => mult_42_n342, A2 => mult_42_n341, B1
                           => mult_42_n343, B2 => mult_42_n320, ZN => 
                           mult_42_n156);
   mult_42_U271 : OAI22_X1 port map( A1 => mult_42_n340, A2 => mult_42_n341, B1
                           => mult_42_n342, B2 => mult_42_n320, ZN => 
                           mult_42_n157);
   mult_42_U270 : OAI22_X1 port map( A1 => mult_42_n336, A2 => mult_42_n337, B1
                           => mult_42_n338, B2 => mult_42_n339, ZN => 
                           mult_42_n19);
   mult_42_U269 : OAI22_X1 port map( A1 => mult_42_n334, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n335, ZN => 
                           mult_42_n25);
   mult_42_U268 : OAI22_X1 port map( A1 => mult_42_n330, A2 => mult_42_n331, B1
                           => mult_42_n332, B2 => mult_42_n333, ZN => 
                           mult_42_n35);
   mult_42_U267 : XOR2_X1 port map( A => B(8), B => x_vector_3_port, Z => 
                           mult_42_n323);
   mult_42_U266 : AOI22_X1 port map( A1 => mult_42_n323, A2 => mult_42_n318, B1
                           => mult_42_n319, B2 => mult_42_n329, ZN => 
                           mult_42_n50);
   mult_42_U265 : OAI22_X1 port map( A1 => mult_42_n325, A2 => mult_42_n326, B1
                           => mult_42_n327, B2 => mult_42_n328, ZN => 
                           mult_42_n321);
   mult_42_U264 : AOI22_X1 port map( A1 => mult_42_n306, A2 => mult_42_n318, B1
                           => mult_42_n319, B2 => mult_42_n323, ZN => 
                           mult_42_n322);
   mult_42_U263 : NAND2_X1 port map( A1 => mult_42_n310, A2 => mult_42_n322, ZN
                           => mult_42_n57);
   mult_42_U262 : XOR2_X1 port map( A => mult_42_n321, B => mult_42_n322, Z => 
                           mult_42_n58);
   mult_42_U261 : XNOR2_X2 port map( A => x_vector_8_port, B => x_vector_7_port
                           , ZN => mult_42_n338);
   mult_42_U260 : XNOR2_X2 port map( A => x_vector_6_port, B => x_vector_5_port
                           , ZN => mult_42_n327);
   mult_42_U259 : XNOR2_X2 port map( A => x_vector_4_port, B => x_vector_3_port
                           , ZN => mult_42_n332);
   mult_42_U258 : INV_X1 port map( A => B(1), ZN => mult_42_n312);
   mult_42_U257 : INV_X1 port map( A => B(0), ZN => mult_42_n313);
   mult_42_U256 : INV_X1 port map( A => x_vector_3_port, ZN => mult_42_n317);
   mult_42_U255 : INV_X1 port map( A => x_vector_0_port, ZN => mult_42_n320);
   mult_42_U254 : INV_X1 port map( A => x_vector_7_port, ZN => mult_42_n315);
   mult_42_U253 : INV_X1 port map( A => x_vector_5_port, ZN => mult_42_n316);
   mult_42_U252 : INV_X1 port map( A => x_vector_9_port, ZN => mult_42_n314);
   mult_42_U251 : INV_X1 port map( A => mult_42_n374, ZN => mult_42_n300);
   mult_42_U250 : INV_X1 port map( A => mult_42_n25, ZN => mult_42_n301);
   mult_42_U249 : INV_X1 port map( A => mult_42_n90, ZN => mult_42_n311);
   mult_42_U248 : INV_X1 port map( A => mult_42_n50, ZN => mult_42_n297);
   mult_42_U247 : INV_X1 port map( A => mult_42_n367, ZN => mult_42_n298);
   mult_42_U246 : INV_X1 port map( A => mult_42_n349, ZN => mult_42_n295);
   mult_42_U245 : INV_X1 port map( A => mult_42_n383, ZN => mult_42_n302);
   mult_42_U244 : INV_X1 port map( A => mult_42_n35, ZN => mult_42_n299);
   mult_42_U243 : INV_X1 port map( A => mult_42_n351, ZN => mult_42_n318);
   mult_42_U242 : INV_X1 port map( A => mult_42_n352, ZN => mult_42_n319);
   mult_42_U241 : INV_X1 port map( A => mult_42_n324, ZN => mult_42_n306);
   mult_42_U240 : INV_X1 port map( A => mult_42_n84, ZN => mult_42_n308);
   mult_42_U239 : INV_X1 port map( A => mult_42_n87, ZN => mult_42_n309);
   mult_42_U238 : INV_X1 port map( A => mult_42_n19, ZN => mult_42_n303);
   mult_42_U237 : INV_X1 port map( A => mult_42_n321, ZN => mult_42_n310);
   mult_42_U236 : INV_X1 port map( A => mult_42_n1, ZN => N12);
   mult_42_U235 : INV_X1 port map( A => mult_42_n74, ZN => mult_42_n305);
   mult_42_U234 : INV_X1 port map( A => mult_42_n79, ZN => mult_42_n307);
   mult_42_U233 : INV_X1 port map( A => mult_42_n60, ZN => mult_42_n296);
   mult_42_U232 : INV_X1 port map( A => mult_42_n67, ZN => mult_42_n304);
   mult_42_U56 : HA_X1 port map( A => mult_42_n148, B => mult_42_n157, CO => 
                           mult_42_n89, S => mult_42_n90);
   mult_42_U55 : FA_X1 port map( A => mult_42_n156, B => mult_42_n139, CI => 
                           mult_42_n147, CO => mult_42_n87, S => mult_42_n88);
   mult_42_U54 : HA_X1 port map( A => mult_42_n107, B => mult_42_n138, CO => 
                           mult_42_n85, S => mult_42_n86);
   mult_42_U53 : FA_X1 port map( A => mult_42_n146, B => mult_42_n155, CI => 
                           mult_42_n86, CO => mult_42_n83, S => mult_42_n84);
   mult_42_U52 : FA_X1 port map( A => mult_42_n154, B => mult_42_n129, CI => 
                           mult_42_n145, CO => mult_42_n81, S => mult_42_n82);
   mult_42_U51 : FA_X1 port map( A => mult_42_n85, B => mult_42_n137, CI => 
                           mult_42_n82, CO => mult_42_n79, S => mult_42_n80);
   mult_42_U50 : HA_X1 port map( A => mult_42_n106, B => mult_42_n128, CO => 
                           mult_42_n77, S => mult_42_n78);
   mult_42_U49 : FA_X1 port map( A => mult_42_n136, B => mult_42_n153, CI => 
                           mult_42_n144, CO => mult_42_n75, S => mult_42_n76);
   mult_42_U48 : FA_X1 port map( A => mult_42_n81, B => mult_42_n78, CI => 
                           mult_42_n76, CO => mult_42_n73, S => mult_42_n74);
   mult_42_U47 : FA_X1 port map( A => mult_42_n135, B => mult_42_n119, CI => 
                           mult_42_n152, CO => mult_42_n71, S => mult_42_n72);
   mult_42_U46 : FA_X1 port map( A => mult_42_n127, B => mult_42_n143, CI => 
                           mult_42_n77, CO => mult_42_n69, S => mult_42_n70);
   mult_42_U45 : FA_X1 port map( A => mult_42_n72, B => mult_42_n75, CI => 
                           mult_42_n70, CO => mult_42_n67, S => mult_42_n68);
   mult_42_U44 : HA_X1 port map( A => mult_42_n105, B => mult_42_n118, CO => 
                           mult_42_n65, S => mult_42_n66);
   mult_42_U43 : FA_X1 port map( A => mult_42_n126, B => mult_42_n134, CI => 
                           mult_42_n142, CO => mult_42_n63, S => mult_42_n64);
   mult_42_U42 : FA_X1 port map( A => mult_42_n66, B => mult_42_n151, CI => 
                           mult_42_n71, CO => mult_42_n61, S => mult_42_n62);
   mult_42_U41 : FA_X1 port map( A => mult_42_n64, B => mult_42_n69, CI => 
                           mult_42_n62, CO => mult_42_n59, S => mult_42_n60);
   mult_42_U38 : FA_X1 port map( A => mult_42_n133, B => mult_42_n117, CI => 
                           mult_42_n295, CO => mult_42_n55, S => mult_42_n56);
   mult_42_U37 : FA_X1 port map( A => mult_42_n58, B => mult_42_n65, CI => 
                           mult_42_n63, CO => mult_42_n53, S => mult_42_n54);
   mult_42_U36 : FA_X1 port map( A => mult_42_n61, B => mult_42_n56, CI => 
                           mult_42_n54, CO => mult_42_n51, S => mult_42_n52);
   mult_42_U34 : FA_X1 port map( A => mult_42_n124, B => mult_42_n116, CI => 
                           mult_42_n132, CO => mult_42_n47, S => mult_42_n48);
   mult_42_U33 : FA_X1 port map( A => mult_42_n57, B => mult_42_n50, CI => 
                           mult_42_n55, CO => mult_42_n45, S => mult_42_n46);
   mult_42_U32 : FA_X1 port map( A => mult_42_n53, B => mult_42_n48, CI => 
                           mult_42_n46, CO => mult_42_n43, S => mult_42_n44);
   mult_42_U31 : FA_X1 port map( A => mult_42_n123, B => mult_42_n115, CI => 
                           mult_42_n140, CO => mult_42_n41, S => mult_42_n42);
   mult_42_U30 : FA_X1 port map( A => mult_42_n297, B => mult_42_n131, CI => 
                           mult_42_n47, CO => mult_42_n39, S => mult_42_n40);
   mult_42_U29 : FA_X1 port map( A => mult_42_n45, B => mult_42_n42, CI => 
                           mult_42_n40, CO => mult_42_n37, S => mult_42_n38);
   mult_42_U27 : FA_X1 port map( A => mult_42_n114, B => mult_42_n122, CI => 
                           mult_42_n299, CO => mult_42_n33, S => mult_42_n34);
   mult_42_U26 : FA_X1 port map( A => mult_42_n34, B => mult_42_n41, CI => 
                           mult_42_n39, CO => mult_42_n31, S => mult_42_n32);
   mult_42_U25 : FA_X1 port map( A => mult_42_n121, B => mult_42_n35, CI => 
                           mult_42_n298, CO => mult_42_n29, S => mult_42_n30);
   mult_42_U24 : FA_X1 port map( A => mult_42_n33, B => mult_42_n113, CI => 
                           mult_42_n30, CO => mult_42_n27, S => mult_42_n28);
   mult_42_U22 : FA_X1 port map( A => mult_42_n301, B => mult_42_n112, CI => 
                           mult_42_n29, CO => mult_42_n23, S => mult_42_n24);
   mult_42_U21 : FA_X1 port map( A => mult_42_n111, B => mult_42_n25, CI => 
                           mult_42_n300, CO => mult_42_n21, S => mult_42_n22);
   mult_42_U10 : FA_X1 port map( A => mult_42_n52, B => mult_42_n59, CI => 
                           mult_42_n10, CO => mult_42_n9, S => N3);
   mult_42_U9 : FA_X1 port map( A => mult_42_n44, B => mult_42_n51, CI => 
                           mult_42_n9, CO => mult_42_n8, S => N4);
   mult_42_U8 : FA_X1 port map( A => mult_42_n38, B => mult_42_n43, CI => 
                           mult_42_n8, CO => mult_42_n7, S => N5);
   mult_42_U7 : FA_X1 port map( A => mult_42_n32, B => mult_42_n37, CI => 
                           mult_42_n7, CO => mult_42_n6, S => N6);
   mult_42_U6 : FA_X1 port map( A => mult_42_n28, B => mult_42_n31, CI => 
                           mult_42_n6, CO => mult_42_n5, S => N7);
   mult_42_U5 : FA_X1 port map( A => mult_42_n24, B => mult_42_n27, CI => 
                           mult_42_n5, CO => mult_42_n4, S => N8);
   mult_42_U4 : FA_X1 port map( A => mult_42_n23, B => mult_42_n22, CI => 
                           mult_42_n4, CO => mult_42_n3, S => N9);
   mult_42_U3 : FA_X1 port map( A => mult_42_n21, B => mult_42_n303, CI => 
                           mult_42_n3, CO => mult_42_n2, S => N10);
   mult_42_U2 : FA_X1 port map( A => mult_42_n302, B => mult_42_n19, CI => 
                           mult_42_n2, CO => mult_42_n1, S => N11);
   mult_42_I2_U391 : NAND2_X1 port map( A1 => x_vector_11_port, A2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n341);
   mult_42_I2_U390 : XNOR2_X1 port map( A => B(12), B => x_vector_11_port, ZN 
                           => mult_42_I2_n340);
   mult_42_I2_U389 : OAI22_X1 port map( A1 => B(11), A2 => mult_42_I2_n341, B1 
                           => mult_42_I2_n340, B2 => mult_42_I2_n320, ZN => 
                           mult_42_I2_n402);
   mult_42_I2_U388 : NAND3_X1 port map( A1 => mult_42_I2_n402, A2 => 
                           mult_42_I2_n312, A3 => x_vector_11_port, ZN => 
                           mult_42_I2_n400);
   mult_42_I2_U387 : XNOR2_X1 port map( A => x_vector_12_port, B => 
                           x_vector_11_port, ZN => mult_42_I2_n352);
   mult_42_I2_U386 : NAND2_X1 port map( A1 => mult_42_I2_n319, A2 => 
                           mult_42_I2_n402, ZN => mult_42_I2_n401);
   mult_42_I2_U385 : MUX2_X1 port map( A => mult_42_I2_n400, B => 
                           mult_42_I2_n401, S => B(10), Z => mult_42_I2_n396);
   mult_42_I2_U384 : XOR2_X1 port map( A => x_vector_13_port, B => 
                           x_vector_12_port, Z => mult_42_I2_n399);
   mult_42_I2_U383 : NAND2_X1 port map( A1 => mult_42_I2_n352, A2 => 
                           mult_42_I2_n399, ZN => mult_42_I2_n351);
   mult_42_I2_U382 : NOR3_X1 port map( A1 => mult_42_I2_n352, A2 => B(10), A3 
                           => mult_42_I2_n317, ZN => mult_42_I2_n398);
   mult_42_I2_U381 : AOI21_X1 port map( B1 => x_vector_13_port, B2 => 
                           mult_42_I2_n318, A => mult_42_I2_n398, ZN => 
                           mult_42_I2_n397);
   mult_42_I2_U380 : OAI222_X1 port map( A1 => mult_42_I2_n396, A2 => 
                           mult_42_I2_n311, B1 => mult_42_I2_n397, B2 => 
                           mult_42_I2_n396, C1 => mult_42_I2_n397, C2 => 
                           mult_42_I2_n311, ZN => mult_42_I2_n395);
   mult_42_I2_U379 : AOI222_X1 port map( A1 => mult_42_I2_n395, A2 => 
                           mult_42_I2_n88, B1 => mult_42_I2_n395, B2 => 
                           mult_42_I2_n89, C1 => mult_42_I2_n89, C2 => 
                           mult_42_I2_n88, ZN => mult_42_I2_n394);
   mult_42_I2_U378 : OAI222_X1 port map( A1 => mult_42_I2_n394, A2 => 
                           mult_42_I2_n308, B1 => mult_42_I2_n394, B2 => 
                           mult_42_I2_n309, C1 => mult_42_I2_n309, C2 => 
                           mult_42_I2_n308, ZN => mult_42_I2_n393);
   mult_42_I2_U377 : AOI222_X1 port map( A1 => mult_42_I2_n393, A2 => 
                           mult_42_I2_n80, B1 => mult_42_I2_n393, B2 => 
                           mult_42_I2_n83, C1 => mult_42_I2_n83, C2 => 
                           mult_42_I2_n80, ZN => mult_42_I2_n392);
   mult_42_I2_U376 : OAI222_X1 port map( A1 => mult_42_I2_n392, A2 => 
                           mult_42_I2_n305, B1 => mult_42_I2_n392, B2 => 
                           mult_42_I2_n307, C1 => mult_42_I2_n307, C2 => 
                           mult_42_I2_n305, ZN => mult_42_I2_n391);
   mult_42_I2_U375 : AOI222_X1 port map( A1 => mult_42_I2_n391, A2 => 
                           mult_42_I2_n68, B1 => mult_42_I2_n391, B2 => 
                           mult_42_I2_n73, C1 => mult_42_I2_n73, C2 => 
                           mult_42_I2_n68, ZN => mult_42_I2_n390);
   mult_42_I2_U374 : OAI222_X1 port map( A1 => mult_42_I2_n390, A2 => 
                           mult_42_I2_n296, B1 => mult_42_I2_n390, B2 => 
                           mult_42_I2_n304, C1 => mult_42_I2_n304, C2 => 
                           mult_42_I2_n296, ZN => mult_42_I2_n10);
   mult_42_I2_U373 : XOR2_X1 port map( A => x_vector_19_port, B => 
                           x_vector_18_port, Z => mult_42_I2_n389);
   mult_42_I2_U372 : NAND2_X1 port map( A1 => mult_42_I2_n338, A2 => 
                           mult_42_I2_n389, ZN => mult_42_I2_n337);
   mult_42_I2_U371 : OR3_X1 port map( A1 => mult_42_I2_n338, A2 => B(10), A3 =>
                           mult_42_I2_n314, ZN => mult_42_I2_n388);
   mult_42_I2_U370 : OAI21_X1 port map( B1 => mult_42_I2_n314, B2 => 
                           mult_42_I2_n337, A => mult_42_I2_n388, ZN => 
                           mult_42_I2_n105);
   mult_42_I2_U369 : XOR2_X1 port map( A => x_vector_17_port, B => 
                           x_vector_16_port, Z => mult_42_I2_n387);
   mult_42_I2_U368 : NAND2_X1 port map( A1 => mult_42_I2_n327, A2 => 
                           mult_42_I2_n387, ZN => mult_42_I2_n326);
   mult_42_I2_U367 : OR3_X1 port map( A1 => mult_42_I2_n327, A2 => B(10), A3 =>
                           mult_42_I2_n315, ZN => mult_42_I2_n386);
   mult_42_I2_U366 : OAI21_X1 port map( B1 => mult_42_I2_n315, B2 => 
                           mult_42_I2_n326, A => mult_42_I2_n386, ZN => 
                           mult_42_I2_n106);
   mult_42_I2_U365 : XOR2_X1 port map( A => x_vector_15_port, B => 
                           x_vector_14_port, Z => mult_42_I2_n385);
   mult_42_I2_U364 : NAND2_X1 port map( A1 => mult_42_I2_n332, A2 => 
                           mult_42_I2_n385, ZN => mult_42_I2_n331);
   mult_42_I2_U363 : OR3_X1 port map( A1 => mult_42_I2_n332, A2 => B(10), A3 =>
                           mult_42_I2_n316, ZN => mult_42_I2_n384);
   mult_42_I2_U362 : OAI21_X1 port map( B1 => mult_42_I2_n316, B2 => 
                           mult_42_I2_n331, A => mult_42_I2_n384, ZN => 
                           mult_42_I2_n107);
   mult_42_I2_U361 : XOR2_X1 port map( A => B(19), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n339);
   mult_42_I2_U360 : OAI22_X1 port map( A1 => mult_42_I2_n339, A2 => 
                           mult_42_I2_n338, B1 => mult_42_I2_n337, B2 => 
                           mult_42_I2_n339, ZN => mult_42_I2_n383);
   mult_42_I2_U359 : XOR2_X1 port map( A => B(17), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n382);
   mult_42_I2_U358 : XOR2_X1 port map( A => B(18), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n336);
   mult_42_I2_U357 : OAI22_X1 port map( A1 => mult_42_I2_n382, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n336, ZN => mult_42_I2_n111);
   mult_42_I2_U356 : XOR2_X1 port map( A => B(16), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n381);
   mult_42_I2_U355 : OAI22_X1 port map( A1 => mult_42_I2_n381, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n382, ZN => mult_42_I2_n112);
   mult_42_I2_U354 : XOR2_X1 port map( A => B(15), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n380);
   mult_42_I2_U353 : OAI22_X1 port map( A1 => mult_42_I2_n380, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n381, ZN => mult_42_I2_n113);
   mult_42_I2_U352 : XOR2_X1 port map( A => B(14), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n379);
   mult_42_I2_U351 : OAI22_X1 port map( A1 => mult_42_I2_n379, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n380, ZN => mult_42_I2_n114);
   mult_42_I2_U350 : XOR2_X1 port map( A => B(13), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n378);
   mult_42_I2_U349 : OAI22_X1 port map( A1 => mult_42_I2_n378, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n379, ZN => mult_42_I2_n115);
   mult_42_I2_U348 : XOR2_X1 port map( A => B(12), B => mult_42_I2_n314, Z => 
                           mult_42_I2_n377);
   mult_42_I2_U347 : OAI22_X1 port map( A1 => mult_42_I2_n377, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n378, ZN => mult_42_I2_n116);
   mult_42_I2_U346 : XOR2_X1 port map( A => mult_42_I2_n312, B => 
                           x_vector_19_port, Z => mult_42_I2_n376);
   mult_42_I2_U345 : OAI22_X1 port map( A1 => mult_42_I2_n376, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n377, ZN => mult_42_I2_n117);
   mult_42_I2_U344 : XOR2_X1 port map( A => mult_42_I2_n314, B => B(10), Z => 
                           mult_42_I2_n375);
   mult_42_I2_U343 : OAI22_X1 port map( A1 => mult_42_I2_n375, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n376, ZN => mult_42_I2_n118);
   mult_42_I2_U342 : NOR2_X1 port map( A1 => mult_42_I2_n338, A2 => 
                           mult_42_I2_n313, ZN => mult_42_I2_n119);
   mult_42_I2_U341 : XOR2_X1 port map( A => B(19), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n335);
   mult_42_I2_U340 : OAI22_X1 port map( A1 => mult_42_I2_n335, A2 => 
                           mult_42_I2_n327, B1 => mult_42_I2_n326, B2 => 
                           mult_42_I2_n335, ZN => mult_42_I2_n374);
   mult_42_I2_U339 : XOR2_X1 port map( A => B(17), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n373);
   mult_42_I2_U338 : XOR2_X1 port map( A => B(18), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n334);
   mult_42_I2_U337 : OAI22_X1 port map( A1 => mult_42_I2_n373, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n334, ZN => mult_42_I2_n121);
   mult_42_I2_U336 : XOR2_X1 port map( A => B(16), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n372);
   mult_42_I2_U335 : OAI22_X1 port map( A1 => mult_42_I2_n372, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n373, ZN => mult_42_I2_n122);
   mult_42_I2_U334 : XOR2_X1 port map( A => B(15), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n371);
   mult_42_I2_U333 : OAI22_X1 port map( A1 => mult_42_I2_n371, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n372, ZN => mult_42_I2_n123);
   mult_42_I2_U332 : XOR2_X1 port map( A => B(14), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n328);
   mult_42_I2_U331 : OAI22_X1 port map( A1 => mult_42_I2_n328, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n371, ZN => mult_42_I2_n124);
   mult_42_I2_U330 : XOR2_X1 port map( A => B(12), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n370);
   mult_42_I2_U329 : XOR2_X1 port map( A => B(13), B => mult_42_I2_n315, Z => 
                           mult_42_I2_n325);
   mult_42_I2_U328 : OAI22_X1 port map( A1 => mult_42_I2_n370, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n325, ZN => mult_42_I2_n126);
   mult_42_I2_U327 : XOR2_X1 port map( A => mult_42_I2_n312, B => 
                           x_vector_17_port, Z => mult_42_I2_n369);
   mult_42_I2_U326 : OAI22_X1 port map( A1 => mult_42_I2_n369, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n370, ZN => mult_42_I2_n127);
   mult_42_I2_U325 : XOR2_X1 port map( A => mult_42_I2_n313, B => 
                           x_vector_17_port, Z => mult_42_I2_n368);
   mult_42_I2_U324 : OAI22_X1 port map( A1 => mult_42_I2_n368, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n369, ZN => mult_42_I2_n128);
   mult_42_I2_U323 : NOR2_X1 port map( A1 => mult_42_I2_n327, A2 => 
                           mult_42_I2_n313, ZN => mult_42_I2_n129);
   mult_42_I2_U322 : XOR2_X1 port map( A => B(19), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n333);
   mult_42_I2_U321 : OAI22_X1 port map( A1 => mult_42_I2_n333, A2 => 
                           mult_42_I2_n332, B1 => mult_42_I2_n331, B2 => 
                           mult_42_I2_n333, ZN => mult_42_I2_n367);
   mult_42_I2_U320 : XOR2_X1 port map( A => B(17), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n366);
   mult_42_I2_U319 : XOR2_X1 port map( A => B(18), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n330);
   mult_42_I2_U318 : OAI22_X1 port map( A1 => mult_42_I2_n366, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n330, ZN => mult_42_I2_n131);
   mult_42_I2_U317 : XOR2_X1 port map( A => B(16), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n365);
   mult_42_I2_U316 : OAI22_X1 port map( A1 => mult_42_I2_n365, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n366, ZN => mult_42_I2_n132);
   mult_42_I2_U315 : XOR2_X1 port map( A => B(15), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n364);
   mult_42_I2_U314 : OAI22_X1 port map( A1 => mult_42_I2_n364, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n365, ZN => mult_42_I2_n133);
   mult_42_I2_U313 : XOR2_X1 port map( A => B(14), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n363);
   mult_42_I2_U312 : OAI22_X1 port map( A1 => mult_42_I2_n363, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n364, ZN => mult_42_I2_n134);
   mult_42_I2_U311 : XOR2_X1 port map( A => B(13), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n362);
   mult_42_I2_U310 : OAI22_X1 port map( A1 => mult_42_I2_n362, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n363, ZN => mult_42_I2_n135);
   mult_42_I2_U309 : XOR2_X1 port map( A => B(12), B => mult_42_I2_n316, Z => 
                           mult_42_I2_n361);
   mult_42_I2_U308 : OAI22_X1 port map( A1 => mult_42_I2_n361, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n362, ZN => mult_42_I2_n136);
   mult_42_I2_U307 : XOR2_X1 port map( A => mult_42_I2_n312, B => 
                           x_vector_15_port, Z => mult_42_I2_n360);
   mult_42_I2_U306 : OAI22_X1 port map( A1 => mult_42_I2_n360, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n361, ZN => mult_42_I2_n137);
   mult_42_I2_U305 : XOR2_X1 port map( A => mult_42_I2_n313, B => 
                           x_vector_15_port, Z => mult_42_I2_n359);
   mult_42_I2_U304 : OAI22_X1 port map( A1 => mult_42_I2_n359, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n360, ZN => mult_42_I2_n138);
   mult_42_I2_U303 : NOR2_X1 port map( A1 => mult_42_I2_n332, A2 => 
                           mult_42_I2_n313, ZN => mult_42_I2_n139);
   mult_42_I2_U302 : XOR2_X1 port map( A => B(19), B => x_vector_13_port, Z => 
                           mult_42_I2_n329);
   mult_42_I2_U301 : AOI22_X1 port map( A1 => mult_42_I2_n329, A2 => 
                           mult_42_I2_n319, B1 => mult_42_I2_n318, B2 => 
                           mult_42_I2_n329, ZN => mult_42_I2_n140);
   mult_42_I2_U300 : XOR2_X1 port map( A => B(16), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n358);
   mult_42_I2_U299 : XOR2_X1 port map( A => B(17), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n324);
   mult_42_I2_U298 : OAI22_X1 port map( A1 => mult_42_I2_n358, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n324, ZN => mult_42_I2_n142);
   mult_42_I2_U297 : XOR2_X1 port map( A => B(15), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n357);
   mult_42_I2_U296 : OAI22_X1 port map( A1 => mult_42_I2_n357, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n358, ZN => mult_42_I2_n143);
   mult_42_I2_U295 : XOR2_X1 port map( A => B(14), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n356);
   mult_42_I2_U294 : OAI22_X1 port map( A1 => mult_42_I2_n356, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n357, ZN => mult_42_I2_n144);
   mult_42_I2_U293 : XOR2_X1 port map( A => B(13), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n355);
   mult_42_I2_U292 : OAI22_X1 port map( A1 => mult_42_I2_n355, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n356, ZN => mult_42_I2_n145);
   mult_42_I2_U291 : XOR2_X1 port map( A => B(12), B => mult_42_I2_n317, Z => 
                           mult_42_I2_n354);
   mult_42_I2_U290 : OAI22_X1 port map( A1 => mult_42_I2_n354, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n355, ZN => mult_42_I2_n146);
   mult_42_I2_U289 : XOR2_X1 port map( A => mult_42_I2_n312, B => 
                           x_vector_13_port, Z => mult_42_I2_n353);
   mult_42_I2_U288 : OAI22_X1 port map( A1 => mult_42_I2_n353, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n354, ZN => mult_42_I2_n147);
   mult_42_I2_U287 : XOR2_X1 port map( A => mult_42_I2_n313, B => 
                           x_vector_13_port, Z => mult_42_I2_n350);
   mult_42_I2_U286 : OAI22_X1 port map( A1 => mult_42_I2_n350, A2 => 
                           mult_42_I2_n351, B1 => mult_42_I2_n352, B2 => 
                           mult_42_I2_n353, ZN => mult_42_I2_n148);
   mult_42_I2_U285 : XNOR2_X1 port map( A => B(19), B => x_vector_11_port, ZN 
                           => mult_42_I2_n348);
   mult_42_I2_U284 : OAI22_X1 port map( A1 => mult_42_I2_n320, A2 => 
                           mult_42_I2_n348, B1 => mult_42_I2_n341, B2 => 
                           mult_42_I2_n348, ZN => mult_42_I2_n349);
   mult_42_I2_U283 : XNOR2_X1 port map( A => B(18), B => x_vector_11_port, ZN 
                           => mult_42_I2_n347);
   mult_42_I2_U282 : OAI22_X1 port map( A1 => mult_42_I2_n347, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n348, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n151);
   mult_42_I2_U281 : XNOR2_X1 port map( A => B(17), B => x_vector_11_port, ZN 
                           => mult_42_I2_n346);
   mult_42_I2_U280 : OAI22_X1 port map( A1 => mult_42_I2_n346, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n347, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n152);
   mult_42_I2_U279 : XNOR2_X1 port map( A => B(16), B => x_vector_11_port, ZN 
                           => mult_42_I2_n345);
   mult_42_I2_U278 : OAI22_X1 port map( A1 => mult_42_I2_n345, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n346, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n153);
   mult_42_I2_U277 : XNOR2_X1 port map( A => B(15), B => x_vector_11_port, ZN 
                           => mult_42_I2_n344);
   mult_42_I2_U276 : OAI22_X1 port map( A1 => mult_42_I2_n344, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n345, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n154);
   mult_42_I2_U275 : XNOR2_X1 port map( A => B(14), B => x_vector_11_port, ZN 
                           => mult_42_I2_n343);
   mult_42_I2_U274 : OAI22_X1 port map( A1 => mult_42_I2_n343, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n344, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n155);
   mult_42_I2_U273 : XNOR2_X1 port map( A => B(13), B => x_vector_11_port, ZN 
                           => mult_42_I2_n342);
   mult_42_I2_U272 : OAI22_X1 port map( A1 => mult_42_I2_n342, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n343, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n156);
   mult_42_I2_U271 : OAI22_X1 port map( A1 => mult_42_I2_n340, A2 => 
                           mult_42_I2_n341, B1 => mult_42_I2_n342, B2 => 
                           mult_42_I2_n320, ZN => mult_42_I2_n157);
   mult_42_I2_U270 : OAI22_X1 port map( A1 => mult_42_I2_n336, A2 => 
                           mult_42_I2_n337, B1 => mult_42_I2_n338, B2 => 
                           mult_42_I2_n339, ZN => mult_42_I2_n19);
   mult_42_I2_U269 : OAI22_X1 port map( A1 => mult_42_I2_n334, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n335, ZN => mult_42_I2_n25);
   mult_42_I2_U268 : OAI22_X1 port map( A1 => mult_42_I2_n330, A2 => 
                           mult_42_I2_n331, B1 => mult_42_I2_n332, B2 => 
                           mult_42_I2_n333, ZN => mult_42_I2_n35);
   mult_42_I2_U267 : XOR2_X1 port map( A => B(18), B => x_vector_13_port, Z => 
                           mult_42_I2_n323);
   mult_42_I2_U266 : AOI22_X1 port map( A1 => mult_42_I2_n323, A2 => 
                           mult_42_I2_n318, B1 => mult_42_I2_n319, B2 => 
                           mult_42_I2_n329, ZN => mult_42_I2_n50);
   mult_42_I2_U265 : OAI22_X1 port map( A1 => mult_42_I2_n325, A2 => 
                           mult_42_I2_n326, B1 => mult_42_I2_n327, B2 => 
                           mult_42_I2_n328, ZN => mult_42_I2_n321);
   mult_42_I2_U264 : AOI22_X1 port map( A1 => mult_42_I2_n306, A2 => 
                           mult_42_I2_n318, B1 => mult_42_I2_n319, B2 => 
                           mult_42_I2_n323, ZN => mult_42_I2_n322);
   mult_42_I2_U263 : NAND2_X1 port map( A1 => mult_42_I2_n310, A2 => 
                           mult_42_I2_n322, ZN => mult_42_I2_n57);
   mult_42_I2_U262 : XOR2_X1 port map( A => mult_42_I2_n321, B => 
                           mult_42_I2_n322, Z => mult_42_I2_n58);
   mult_42_I2_U261 : XNOR2_X2 port map( A => x_vector_18_port, B => 
                           x_vector_17_port, ZN => mult_42_I2_n338);
   mult_42_I2_U260 : XNOR2_X2 port map( A => x_vector_16_port, B => 
                           x_vector_15_port, ZN => mult_42_I2_n327);
   mult_42_I2_U259 : XNOR2_X2 port map( A => x_vector_14_port, B => 
                           x_vector_13_port, ZN => mult_42_I2_n332);
   mult_42_I2_U258 : INV_X1 port map( A => B(11), ZN => mult_42_I2_n312);
   mult_42_I2_U257 : INV_X1 port map( A => B(10), ZN => mult_42_I2_n313);
   mult_42_I2_U256 : INV_X1 port map( A => x_vector_13_port, ZN => 
                           mult_42_I2_n317);
   mult_42_I2_U255 : INV_X1 port map( A => x_vector_10_port, ZN => 
                           mult_42_I2_n320);
   mult_42_I2_U254 : INV_X1 port map( A => x_vector_17_port, ZN => 
                           mult_42_I2_n315);
   mult_42_I2_U253 : INV_X1 port map( A => x_vector_15_port, ZN => 
                           mult_42_I2_n316);
   mult_42_I2_U252 : INV_X1 port map( A => x_vector_19_port, ZN => 
                           mult_42_I2_n314);
   mult_42_I2_U251 : INV_X1 port map( A => mult_42_I2_n374, ZN => 
                           mult_42_I2_n300);
   mult_42_I2_U250 : INV_X1 port map( A => mult_42_I2_n25, ZN => 
                           mult_42_I2_n301);
   mult_42_I2_U249 : INV_X1 port map( A => mult_42_I2_n90, ZN => 
                           mult_42_I2_n311);
   mult_42_I2_U248 : INV_X1 port map( A => mult_42_I2_n50, ZN => 
                           mult_42_I2_n297);
   mult_42_I2_U247 : INV_X1 port map( A => mult_42_I2_n367, ZN => 
                           mult_42_I2_n298);
   mult_42_I2_U246 : INV_X1 port map( A => mult_42_I2_n349, ZN => 
                           mult_42_I2_n295);
   mult_42_I2_U245 : INV_X1 port map( A => mult_42_I2_n383, ZN => 
                           mult_42_I2_n302);
   mult_42_I2_U244 : INV_X1 port map( A => mult_42_I2_n35, ZN => 
                           mult_42_I2_n299);
   mult_42_I2_U243 : INV_X1 port map( A => mult_42_I2_n351, ZN => 
                           mult_42_I2_n318);
   mult_42_I2_U242 : INV_X1 port map( A => mult_42_I2_n352, ZN => 
                           mult_42_I2_n319);
   mult_42_I2_U241 : INV_X1 port map( A => mult_42_I2_n324, ZN => 
                           mult_42_I2_n306);
   mult_42_I2_U240 : INV_X1 port map( A => mult_42_I2_n84, ZN => 
                           mult_42_I2_n308);
   mult_42_I2_U239 : INV_X1 port map( A => mult_42_I2_n87, ZN => 
                           mult_42_I2_n309);
   mult_42_I2_U238 : INV_X1 port map( A => mult_42_I2_n19, ZN => 
                           mult_42_I2_n303);
   mult_42_I2_U237 : INV_X1 port map( A => mult_42_I2_n321, ZN => 
                           mult_42_I2_n310);
   mult_42_I2_U236 : INV_X1 port map( A => mult_42_I2_n1, ZN => N22);
   mult_42_I2_U235 : INV_X1 port map( A => mult_42_I2_n74, ZN => 
                           mult_42_I2_n305);
   mult_42_I2_U234 : INV_X1 port map( A => mult_42_I2_n79, ZN => 
                           mult_42_I2_n307);
   mult_42_I2_U233 : INV_X1 port map( A => mult_42_I2_n60, ZN => 
                           mult_42_I2_n296);
   mult_42_I2_U232 : INV_X1 port map( A => mult_42_I2_n67, ZN => 
                           mult_42_I2_n304);
   mult_42_I2_U56 : HA_X1 port map( A => mult_42_I2_n148, B => mult_42_I2_n157,
                           CO => mult_42_I2_n89, S => mult_42_I2_n90);
   mult_42_I2_U55 : FA_X1 port map( A => mult_42_I2_n156, B => mult_42_I2_n139,
                           CI => mult_42_I2_n147, CO => mult_42_I2_n87, S => 
                           mult_42_I2_n88);
   mult_42_I2_U54 : HA_X1 port map( A => mult_42_I2_n107, B => mult_42_I2_n138,
                           CO => mult_42_I2_n85, S => mult_42_I2_n86);
   mult_42_I2_U53 : FA_X1 port map( A => mult_42_I2_n146, B => mult_42_I2_n155,
                           CI => mult_42_I2_n86, CO => mult_42_I2_n83, S => 
                           mult_42_I2_n84);
   mult_42_I2_U52 : FA_X1 port map( A => mult_42_I2_n154, B => mult_42_I2_n129,
                           CI => mult_42_I2_n145, CO => mult_42_I2_n81, S => 
                           mult_42_I2_n82);
   mult_42_I2_U51 : FA_X1 port map( A => mult_42_I2_n85, B => mult_42_I2_n137, 
                           CI => mult_42_I2_n82, CO => mult_42_I2_n79, S => 
                           mult_42_I2_n80);
   mult_42_I2_U50 : HA_X1 port map( A => mult_42_I2_n106, B => mult_42_I2_n128,
                           CO => mult_42_I2_n77, S => mult_42_I2_n78);
   mult_42_I2_U49 : FA_X1 port map( A => mult_42_I2_n136, B => mult_42_I2_n153,
                           CI => mult_42_I2_n144, CO => mult_42_I2_n75, S => 
                           mult_42_I2_n76);
   mult_42_I2_U48 : FA_X1 port map( A => mult_42_I2_n81, B => mult_42_I2_n78, 
                           CI => mult_42_I2_n76, CO => mult_42_I2_n73, S => 
                           mult_42_I2_n74);
   mult_42_I2_U47 : FA_X1 port map( A => mult_42_I2_n135, B => mult_42_I2_n119,
                           CI => mult_42_I2_n152, CO => mult_42_I2_n71, S => 
                           mult_42_I2_n72);
   mult_42_I2_U46 : FA_X1 port map( A => mult_42_I2_n127, B => mult_42_I2_n143,
                           CI => mult_42_I2_n77, CO => mult_42_I2_n69, S => 
                           mult_42_I2_n70);
   mult_42_I2_U45 : FA_X1 port map( A => mult_42_I2_n72, B => mult_42_I2_n75, 
                           CI => mult_42_I2_n70, CO => mult_42_I2_n67, S => 
                           mult_42_I2_n68);
   mult_42_I2_U44 : HA_X1 port map( A => mult_42_I2_n105, B => mult_42_I2_n118,
                           CO => mult_42_I2_n65, S => mult_42_I2_n66);
   mult_42_I2_U43 : FA_X1 port map( A => mult_42_I2_n126, B => mult_42_I2_n134,
                           CI => mult_42_I2_n142, CO => mult_42_I2_n63, S => 
                           mult_42_I2_n64);
   mult_42_I2_U42 : FA_X1 port map( A => mult_42_I2_n66, B => mult_42_I2_n151, 
                           CI => mult_42_I2_n71, CO => mult_42_I2_n61, S => 
                           mult_42_I2_n62);
   mult_42_I2_U41 : FA_X1 port map( A => mult_42_I2_n64, B => mult_42_I2_n69, 
                           CI => mult_42_I2_n62, CO => mult_42_I2_n59, S => 
                           mult_42_I2_n60);
   mult_42_I2_U38 : FA_X1 port map( A => mult_42_I2_n133, B => mult_42_I2_n117,
                           CI => mult_42_I2_n295, CO => mult_42_I2_n55, S => 
                           mult_42_I2_n56);
   mult_42_I2_U37 : FA_X1 port map( A => mult_42_I2_n58, B => mult_42_I2_n65, 
                           CI => mult_42_I2_n63, CO => mult_42_I2_n53, S => 
                           mult_42_I2_n54);
   mult_42_I2_U36 : FA_X1 port map( A => mult_42_I2_n61, B => mult_42_I2_n56, 
                           CI => mult_42_I2_n54, CO => mult_42_I2_n51, S => 
                           mult_42_I2_n52);
   mult_42_I2_U34 : FA_X1 port map( A => mult_42_I2_n124, B => mult_42_I2_n116,
                           CI => mult_42_I2_n132, CO => mult_42_I2_n47, S => 
                           mult_42_I2_n48);
   mult_42_I2_U33 : FA_X1 port map( A => mult_42_I2_n57, B => mult_42_I2_n50, 
                           CI => mult_42_I2_n55, CO => mult_42_I2_n45, S => 
                           mult_42_I2_n46);
   mult_42_I2_U32 : FA_X1 port map( A => mult_42_I2_n53, B => mult_42_I2_n48, 
                           CI => mult_42_I2_n46, CO => mult_42_I2_n43, S => 
                           mult_42_I2_n44);
   mult_42_I2_U31 : FA_X1 port map( A => mult_42_I2_n123, B => mult_42_I2_n115,
                           CI => mult_42_I2_n140, CO => mult_42_I2_n41, S => 
                           mult_42_I2_n42);
   mult_42_I2_U30 : FA_X1 port map( A => mult_42_I2_n297, B => mult_42_I2_n131,
                           CI => mult_42_I2_n47, CO => mult_42_I2_n39, S => 
                           mult_42_I2_n40);
   mult_42_I2_U29 : FA_X1 port map( A => mult_42_I2_n45, B => mult_42_I2_n42, 
                           CI => mult_42_I2_n40, CO => mult_42_I2_n37, S => 
                           mult_42_I2_n38);
   mult_42_I2_U27 : FA_X1 port map( A => mult_42_I2_n114, B => mult_42_I2_n122,
                           CI => mult_42_I2_n299, CO => mult_42_I2_n33, S => 
                           mult_42_I2_n34);
   mult_42_I2_U26 : FA_X1 port map( A => mult_42_I2_n34, B => mult_42_I2_n41, 
                           CI => mult_42_I2_n39, CO => mult_42_I2_n31, S => 
                           mult_42_I2_n32);
   mult_42_I2_U25 : FA_X1 port map( A => mult_42_I2_n121, B => mult_42_I2_n35, 
                           CI => mult_42_I2_n298, CO => mult_42_I2_n29, S => 
                           mult_42_I2_n30);
   mult_42_I2_U24 : FA_X1 port map( A => mult_42_I2_n33, B => mult_42_I2_n113, 
                           CI => mult_42_I2_n30, CO => mult_42_I2_n27, S => 
                           mult_42_I2_n28);
   mult_42_I2_U22 : FA_X1 port map( A => mult_42_I2_n301, B => mult_42_I2_n112,
                           CI => mult_42_I2_n29, CO => mult_42_I2_n23, S => 
                           mult_42_I2_n24);
   mult_42_I2_U21 : FA_X1 port map( A => mult_42_I2_n111, B => mult_42_I2_n25, 
                           CI => mult_42_I2_n300, CO => mult_42_I2_n21, S => 
                           mult_42_I2_n22);
   mult_42_I2_U10 : FA_X1 port map( A => mult_42_I2_n52, B => mult_42_I2_n59, 
                           CI => mult_42_I2_n10, CO => mult_42_I2_n9, S => N13)
                           ;
   mult_42_I2_U9 : FA_X1 port map( A => mult_42_I2_n44, B => mult_42_I2_n51, CI
                           => mult_42_I2_n9, CO => mult_42_I2_n8, S => N14);
   mult_42_I2_U8 : FA_X1 port map( A => mult_42_I2_n38, B => mult_42_I2_n43, CI
                           => mult_42_I2_n8, CO => mult_42_I2_n7, S => N15);
   mult_42_I2_U7 : FA_X1 port map( A => mult_42_I2_n32, B => mult_42_I2_n37, CI
                           => mult_42_I2_n7, CO => mult_42_I2_n6, S => N16);
   mult_42_I2_U6 : FA_X1 port map( A => mult_42_I2_n28, B => mult_42_I2_n31, CI
                           => mult_42_I2_n6, CO => mult_42_I2_n5, S => N17);
   mult_42_I2_U5 : FA_X1 port map( A => mult_42_I2_n24, B => mult_42_I2_n27, CI
                           => mult_42_I2_n5, CO => mult_42_I2_n4, S => N18);
   mult_42_I2_U4 : FA_X1 port map( A => mult_42_I2_n23, B => mult_42_I2_n22, CI
                           => mult_42_I2_n4, CO => mult_42_I2_n3, S => N19);
   mult_42_I2_U3 : FA_X1 port map( A => mult_42_I2_n21, B => mult_42_I2_n303, 
                           CI => mult_42_I2_n3, CO => mult_42_I2_n2, S => N20);
   mult_42_I2_U2 : FA_X1 port map( A => mult_42_I2_n302, B => mult_42_I2_n19, 
                           CI => mult_42_I2_n2, CO => mult_42_I2_n1, S => 
                           N21_port);
   mult_42_I3_U391 : NAND2_X1 port map( A1 => x_vector_21_port, A2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n341);
   mult_42_I3_U390 : XNOR2_X1 port map( A => B(22), B => x_vector_21_port, ZN 
                           => mult_42_I3_n340);
   mult_42_I3_U389 : OAI22_X1 port map( A1 => B(21), A2 => mult_42_I3_n341, B1 
                           => mult_42_I3_n340, B2 => mult_42_I3_n320, ZN => 
                           mult_42_I3_n402);
   mult_42_I3_U388 : NAND3_X1 port map( A1 => mult_42_I3_n402, A2 => 
                           mult_42_I3_n312, A3 => x_vector_21_port, ZN => 
                           mult_42_I3_n400);
   mult_42_I3_U387 : XNOR2_X1 port map( A => x_vector_22_port, B => 
                           x_vector_21_port, ZN => mult_42_I3_n352);
   mult_42_I3_U386 : NAND2_X1 port map( A1 => mult_42_I3_n319, A2 => 
                           mult_42_I3_n402, ZN => mult_42_I3_n401);
   mult_42_I3_U385 : MUX2_X1 port map( A => mult_42_I3_n400, B => 
                           mult_42_I3_n401, S => B(20), Z => mult_42_I3_n396);
   mult_42_I3_U384 : XOR2_X1 port map( A => x_vector_23_port, B => 
                           x_vector_22_port, Z => mult_42_I3_n399);
   mult_42_I3_U383 : NAND2_X1 port map( A1 => mult_42_I3_n352, A2 => 
                           mult_42_I3_n399, ZN => mult_42_I3_n351);
   mult_42_I3_U382 : NOR3_X1 port map( A1 => mult_42_I3_n352, A2 => B(20), A3 
                           => mult_42_I3_n317, ZN => mult_42_I3_n398);
   mult_42_I3_U381 : AOI21_X1 port map( B1 => x_vector_23_port, B2 => 
                           mult_42_I3_n318, A => mult_42_I3_n398, ZN => 
                           mult_42_I3_n397);
   mult_42_I3_U380 : OAI222_X1 port map( A1 => mult_42_I3_n396, A2 => 
                           mult_42_I3_n311, B1 => mult_42_I3_n397, B2 => 
                           mult_42_I3_n396, C1 => mult_42_I3_n397, C2 => 
                           mult_42_I3_n311, ZN => mult_42_I3_n395);
   mult_42_I3_U379 : AOI222_X1 port map( A1 => mult_42_I3_n395, A2 => 
                           mult_42_I3_n88, B1 => mult_42_I3_n395, B2 => 
                           mult_42_I3_n89, C1 => mult_42_I3_n89, C2 => 
                           mult_42_I3_n88, ZN => mult_42_I3_n394);
   mult_42_I3_U378 : OAI222_X1 port map( A1 => mult_42_I3_n394, A2 => 
                           mult_42_I3_n308, B1 => mult_42_I3_n394, B2 => 
                           mult_42_I3_n309, C1 => mult_42_I3_n309, C2 => 
                           mult_42_I3_n308, ZN => mult_42_I3_n393);
   mult_42_I3_U377 : AOI222_X1 port map( A1 => mult_42_I3_n393, A2 => 
                           mult_42_I3_n80, B1 => mult_42_I3_n393, B2 => 
                           mult_42_I3_n83, C1 => mult_42_I3_n83, C2 => 
                           mult_42_I3_n80, ZN => mult_42_I3_n392);
   mult_42_I3_U376 : OAI222_X1 port map( A1 => mult_42_I3_n392, A2 => 
                           mult_42_I3_n305, B1 => mult_42_I3_n392, B2 => 
                           mult_42_I3_n307, C1 => mult_42_I3_n307, C2 => 
                           mult_42_I3_n305, ZN => mult_42_I3_n391);
   mult_42_I3_U375 : AOI222_X1 port map( A1 => mult_42_I3_n391, A2 => 
                           mult_42_I3_n68, B1 => mult_42_I3_n391, B2 => 
                           mult_42_I3_n73, C1 => mult_42_I3_n73, C2 => 
                           mult_42_I3_n68, ZN => mult_42_I3_n390);
   mult_42_I3_U374 : OAI222_X1 port map( A1 => mult_42_I3_n390, A2 => 
                           mult_42_I3_n296, B1 => mult_42_I3_n390, B2 => 
                           mult_42_I3_n304, C1 => mult_42_I3_n304, C2 => 
                           mult_42_I3_n296, ZN => mult_42_I3_n10);
   mult_42_I3_U373 : XOR2_X1 port map( A => x_vector_29_port, B => 
                           x_vector_28_port, Z => mult_42_I3_n389);
   mult_42_I3_U372 : NAND2_X1 port map( A1 => mult_42_I3_n338, A2 => 
                           mult_42_I3_n389, ZN => mult_42_I3_n337);
   mult_42_I3_U371 : OR3_X1 port map( A1 => mult_42_I3_n338, A2 => B(20), A3 =>
                           mult_42_I3_n314, ZN => mult_42_I3_n388);
   mult_42_I3_U370 : OAI21_X1 port map( B1 => mult_42_I3_n314, B2 => 
                           mult_42_I3_n337, A => mult_42_I3_n388, ZN => 
                           mult_42_I3_n105);
   mult_42_I3_U369 : XOR2_X1 port map( A => x_vector_27_port, B => 
                           x_vector_26_port, Z => mult_42_I3_n387);
   mult_42_I3_U368 : NAND2_X1 port map( A1 => mult_42_I3_n327, A2 => 
                           mult_42_I3_n387, ZN => mult_42_I3_n326);
   mult_42_I3_U367 : OR3_X1 port map( A1 => mult_42_I3_n327, A2 => B(20), A3 =>
                           mult_42_I3_n315, ZN => mult_42_I3_n386);
   mult_42_I3_U366 : OAI21_X1 port map( B1 => mult_42_I3_n315, B2 => 
                           mult_42_I3_n326, A => mult_42_I3_n386, ZN => 
                           mult_42_I3_n106);
   mult_42_I3_U365 : XOR2_X1 port map( A => x_vector_25_port, B => 
                           x_vector_24_port, Z => mult_42_I3_n385);
   mult_42_I3_U364 : NAND2_X1 port map( A1 => mult_42_I3_n332, A2 => 
                           mult_42_I3_n385, ZN => mult_42_I3_n331);
   mult_42_I3_U363 : OR3_X1 port map( A1 => mult_42_I3_n332, A2 => B(20), A3 =>
                           mult_42_I3_n316, ZN => mult_42_I3_n384);
   mult_42_I3_U362 : OAI21_X1 port map( B1 => mult_42_I3_n316, B2 => 
                           mult_42_I3_n331, A => mult_42_I3_n384, ZN => 
                           mult_42_I3_n107);
   mult_42_I3_U361 : XOR2_X1 port map( A => B(29), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n339);
   mult_42_I3_U360 : OAI22_X1 port map( A1 => mult_42_I3_n339, A2 => 
                           mult_42_I3_n338, B1 => mult_42_I3_n337, B2 => 
                           mult_42_I3_n339, ZN => mult_42_I3_n383);
   mult_42_I3_U359 : XOR2_X1 port map( A => B(27), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n382);
   mult_42_I3_U358 : XOR2_X1 port map( A => B(28), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n336);
   mult_42_I3_U357 : OAI22_X1 port map( A1 => mult_42_I3_n382, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n336, ZN => mult_42_I3_n111);
   mult_42_I3_U356 : XOR2_X1 port map( A => B(26), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n381);
   mult_42_I3_U355 : OAI22_X1 port map( A1 => mult_42_I3_n381, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n382, ZN => mult_42_I3_n112);
   mult_42_I3_U354 : XOR2_X1 port map( A => B(25), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n380);
   mult_42_I3_U353 : OAI22_X1 port map( A1 => mult_42_I3_n380, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n381, ZN => mult_42_I3_n113);
   mult_42_I3_U352 : XOR2_X1 port map( A => B(24), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n379);
   mult_42_I3_U351 : OAI22_X1 port map( A1 => mult_42_I3_n379, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n380, ZN => mult_42_I3_n114);
   mult_42_I3_U350 : XOR2_X1 port map( A => B(23), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n378);
   mult_42_I3_U349 : OAI22_X1 port map( A1 => mult_42_I3_n378, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n379, ZN => mult_42_I3_n115);
   mult_42_I3_U348 : XOR2_X1 port map( A => B(22), B => mult_42_I3_n314, Z => 
                           mult_42_I3_n377);
   mult_42_I3_U347 : OAI22_X1 port map( A1 => mult_42_I3_n377, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n378, ZN => mult_42_I3_n116);
   mult_42_I3_U346 : XOR2_X1 port map( A => mult_42_I3_n312, B => 
                           x_vector_29_port, Z => mult_42_I3_n376);
   mult_42_I3_U345 : OAI22_X1 port map( A1 => mult_42_I3_n376, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n377, ZN => mult_42_I3_n117);
   mult_42_I3_U344 : XOR2_X1 port map( A => mult_42_I3_n314, B => B(20), Z => 
                           mult_42_I3_n375);
   mult_42_I3_U343 : OAI22_X1 port map( A1 => mult_42_I3_n375, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n376, ZN => mult_42_I3_n118);
   mult_42_I3_U342 : NOR2_X1 port map( A1 => mult_42_I3_n338, A2 => 
                           mult_42_I3_n313, ZN => mult_42_I3_n119);
   mult_42_I3_U341 : XOR2_X1 port map( A => B(29), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n335);
   mult_42_I3_U340 : OAI22_X1 port map( A1 => mult_42_I3_n335, A2 => 
                           mult_42_I3_n327, B1 => mult_42_I3_n326, B2 => 
                           mult_42_I3_n335, ZN => mult_42_I3_n374);
   mult_42_I3_U339 : XOR2_X1 port map( A => B(27), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n373);
   mult_42_I3_U338 : XOR2_X1 port map( A => B(28), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n334);
   mult_42_I3_U337 : OAI22_X1 port map( A1 => mult_42_I3_n373, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n334, ZN => mult_42_I3_n121);
   mult_42_I3_U336 : XOR2_X1 port map( A => B(26), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n372);
   mult_42_I3_U335 : OAI22_X1 port map( A1 => mult_42_I3_n372, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n373, ZN => mult_42_I3_n122);
   mult_42_I3_U334 : XOR2_X1 port map( A => B(25), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n371);
   mult_42_I3_U333 : OAI22_X1 port map( A1 => mult_42_I3_n371, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n372, ZN => mult_42_I3_n123);
   mult_42_I3_U332 : XOR2_X1 port map( A => B(24), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n328);
   mult_42_I3_U331 : OAI22_X1 port map( A1 => mult_42_I3_n328, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n371, ZN => mult_42_I3_n124);
   mult_42_I3_U330 : XOR2_X1 port map( A => B(22), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n370);
   mult_42_I3_U329 : XOR2_X1 port map( A => B(23), B => mult_42_I3_n315, Z => 
                           mult_42_I3_n325);
   mult_42_I3_U328 : OAI22_X1 port map( A1 => mult_42_I3_n370, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n325, ZN => mult_42_I3_n126);
   mult_42_I3_U327 : XOR2_X1 port map( A => mult_42_I3_n312, B => 
                           x_vector_27_port, Z => mult_42_I3_n369);
   mult_42_I3_U326 : OAI22_X1 port map( A1 => mult_42_I3_n369, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n370, ZN => mult_42_I3_n127);
   mult_42_I3_U325 : XOR2_X1 port map( A => mult_42_I3_n313, B => 
                           x_vector_27_port, Z => mult_42_I3_n368);
   mult_42_I3_U324 : OAI22_X1 port map( A1 => mult_42_I3_n368, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n369, ZN => mult_42_I3_n128);
   mult_42_I3_U323 : NOR2_X1 port map( A1 => mult_42_I3_n327, A2 => 
                           mult_42_I3_n313, ZN => mult_42_I3_n129);
   mult_42_I3_U322 : XOR2_X1 port map( A => B(29), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n333);
   mult_42_I3_U321 : OAI22_X1 port map( A1 => mult_42_I3_n333, A2 => 
                           mult_42_I3_n332, B1 => mult_42_I3_n331, B2 => 
                           mult_42_I3_n333, ZN => mult_42_I3_n367);
   mult_42_I3_U320 : XOR2_X1 port map( A => B(27), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n366);
   mult_42_I3_U319 : XOR2_X1 port map( A => B(28), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n330);
   mult_42_I3_U318 : OAI22_X1 port map( A1 => mult_42_I3_n366, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n330, ZN => mult_42_I3_n131);
   mult_42_I3_U317 : XOR2_X1 port map( A => B(26), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n365);
   mult_42_I3_U316 : OAI22_X1 port map( A1 => mult_42_I3_n365, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n366, ZN => mult_42_I3_n132);
   mult_42_I3_U315 : XOR2_X1 port map( A => B(25), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n364);
   mult_42_I3_U314 : OAI22_X1 port map( A1 => mult_42_I3_n364, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n365, ZN => mult_42_I3_n133);
   mult_42_I3_U313 : XOR2_X1 port map( A => B(24), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n363);
   mult_42_I3_U312 : OAI22_X1 port map( A1 => mult_42_I3_n363, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n364, ZN => mult_42_I3_n134);
   mult_42_I3_U311 : XOR2_X1 port map( A => B(23), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n362);
   mult_42_I3_U310 : OAI22_X1 port map( A1 => mult_42_I3_n362, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n363, ZN => mult_42_I3_n135);
   mult_42_I3_U309 : XOR2_X1 port map( A => B(22), B => mult_42_I3_n316, Z => 
                           mult_42_I3_n361);
   mult_42_I3_U308 : OAI22_X1 port map( A1 => mult_42_I3_n361, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n362, ZN => mult_42_I3_n136);
   mult_42_I3_U307 : XOR2_X1 port map( A => mult_42_I3_n312, B => 
                           x_vector_25_port, Z => mult_42_I3_n360);
   mult_42_I3_U306 : OAI22_X1 port map( A1 => mult_42_I3_n360, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n361, ZN => mult_42_I3_n137);
   mult_42_I3_U305 : XOR2_X1 port map( A => mult_42_I3_n313, B => 
                           x_vector_25_port, Z => mult_42_I3_n359);
   mult_42_I3_U304 : OAI22_X1 port map( A1 => mult_42_I3_n359, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n360, ZN => mult_42_I3_n138);
   mult_42_I3_U303 : NOR2_X1 port map( A1 => mult_42_I3_n332, A2 => 
                           mult_42_I3_n313, ZN => mult_42_I3_n139);
   mult_42_I3_U302 : XOR2_X1 port map( A => B(29), B => x_vector_23_port, Z => 
                           mult_42_I3_n329);
   mult_42_I3_U301 : AOI22_X1 port map( A1 => mult_42_I3_n329, A2 => 
                           mult_42_I3_n319, B1 => mult_42_I3_n318, B2 => 
                           mult_42_I3_n329, ZN => mult_42_I3_n140);
   mult_42_I3_U300 : XOR2_X1 port map( A => B(26), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n358);
   mult_42_I3_U299 : XOR2_X1 port map( A => B(27), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n324);
   mult_42_I3_U298 : OAI22_X1 port map( A1 => mult_42_I3_n358, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n324, ZN => mult_42_I3_n142);
   mult_42_I3_U297 : XOR2_X1 port map( A => B(25), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n357);
   mult_42_I3_U296 : OAI22_X1 port map( A1 => mult_42_I3_n357, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n358, ZN => mult_42_I3_n143);
   mult_42_I3_U295 : XOR2_X1 port map( A => B(24), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n356);
   mult_42_I3_U294 : OAI22_X1 port map( A1 => mult_42_I3_n356, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n357, ZN => mult_42_I3_n144);
   mult_42_I3_U293 : XOR2_X1 port map( A => B(23), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n355);
   mult_42_I3_U292 : OAI22_X1 port map( A1 => mult_42_I3_n355, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n356, ZN => mult_42_I3_n145);
   mult_42_I3_U291 : XOR2_X1 port map( A => B(22), B => mult_42_I3_n317, Z => 
                           mult_42_I3_n354);
   mult_42_I3_U290 : OAI22_X1 port map( A1 => mult_42_I3_n354, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n355, ZN => mult_42_I3_n146);
   mult_42_I3_U289 : XOR2_X1 port map( A => mult_42_I3_n312, B => 
                           x_vector_23_port, Z => mult_42_I3_n353);
   mult_42_I3_U288 : OAI22_X1 port map( A1 => mult_42_I3_n353, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n354, ZN => mult_42_I3_n147);
   mult_42_I3_U287 : XOR2_X1 port map( A => mult_42_I3_n313, B => 
                           x_vector_23_port, Z => mult_42_I3_n350);
   mult_42_I3_U286 : OAI22_X1 port map( A1 => mult_42_I3_n350, A2 => 
                           mult_42_I3_n351, B1 => mult_42_I3_n352, B2 => 
                           mult_42_I3_n353, ZN => mult_42_I3_n148);
   mult_42_I3_U285 : XNOR2_X1 port map( A => B(29), B => x_vector_21_port, ZN 
                           => mult_42_I3_n348);
   mult_42_I3_U284 : OAI22_X1 port map( A1 => mult_42_I3_n320, A2 => 
                           mult_42_I3_n348, B1 => mult_42_I3_n341, B2 => 
                           mult_42_I3_n348, ZN => mult_42_I3_n349);
   mult_42_I3_U283 : XNOR2_X1 port map( A => B(28), B => x_vector_21_port, ZN 
                           => mult_42_I3_n347);
   mult_42_I3_U282 : OAI22_X1 port map( A1 => mult_42_I3_n347, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n348, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n151);
   mult_42_I3_U281 : XNOR2_X1 port map( A => B(27), B => x_vector_21_port, ZN 
                           => mult_42_I3_n346);
   mult_42_I3_U280 : OAI22_X1 port map( A1 => mult_42_I3_n346, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n347, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n152);
   mult_42_I3_U279 : XNOR2_X1 port map( A => B(26), B => x_vector_21_port, ZN 
                           => mult_42_I3_n345);
   mult_42_I3_U278 : OAI22_X1 port map( A1 => mult_42_I3_n345, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n346, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n153);
   mult_42_I3_U277 : XNOR2_X1 port map( A => B(25), B => x_vector_21_port, ZN 
                           => mult_42_I3_n344);
   mult_42_I3_U276 : OAI22_X1 port map( A1 => mult_42_I3_n344, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n345, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n154);
   mult_42_I3_U275 : XNOR2_X1 port map( A => B(24), B => x_vector_21_port, ZN 
                           => mult_42_I3_n343);
   mult_42_I3_U274 : OAI22_X1 port map( A1 => mult_42_I3_n343, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n344, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n155);
   mult_42_I3_U273 : XNOR2_X1 port map( A => B(23), B => x_vector_21_port, ZN 
                           => mult_42_I3_n342);
   mult_42_I3_U272 : OAI22_X1 port map( A1 => mult_42_I3_n342, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n343, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n156);
   mult_42_I3_U271 : OAI22_X1 port map( A1 => mult_42_I3_n340, A2 => 
                           mult_42_I3_n341, B1 => mult_42_I3_n342, B2 => 
                           mult_42_I3_n320, ZN => mult_42_I3_n157);
   mult_42_I3_U270 : OAI22_X1 port map( A1 => mult_42_I3_n336, A2 => 
                           mult_42_I3_n337, B1 => mult_42_I3_n338, B2 => 
                           mult_42_I3_n339, ZN => mult_42_I3_n19);
   mult_42_I3_U269 : OAI22_X1 port map( A1 => mult_42_I3_n334, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n335, ZN => mult_42_I3_n25);
   mult_42_I3_U268 : OAI22_X1 port map( A1 => mult_42_I3_n330, A2 => 
                           mult_42_I3_n331, B1 => mult_42_I3_n332, B2 => 
                           mult_42_I3_n333, ZN => mult_42_I3_n35);
   mult_42_I3_U267 : XOR2_X1 port map( A => B(28), B => x_vector_23_port, Z => 
                           mult_42_I3_n323);
   mult_42_I3_U266 : AOI22_X1 port map( A1 => mult_42_I3_n323, A2 => 
                           mult_42_I3_n318, B1 => mult_42_I3_n319, B2 => 
                           mult_42_I3_n329, ZN => mult_42_I3_n50);
   mult_42_I3_U265 : OAI22_X1 port map( A1 => mult_42_I3_n325, A2 => 
                           mult_42_I3_n326, B1 => mult_42_I3_n327, B2 => 
                           mult_42_I3_n328, ZN => mult_42_I3_n321);
   mult_42_I3_U264 : AOI22_X1 port map( A1 => mult_42_I3_n306, A2 => 
                           mult_42_I3_n318, B1 => mult_42_I3_n319, B2 => 
                           mult_42_I3_n323, ZN => mult_42_I3_n322);
   mult_42_I3_U263 : NAND2_X1 port map( A1 => mult_42_I3_n310, A2 => 
                           mult_42_I3_n322, ZN => mult_42_I3_n57);
   mult_42_I3_U262 : XOR2_X1 port map( A => mult_42_I3_n321, B => 
                           mult_42_I3_n322, Z => mult_42_I3_n58);
   mult_42_I3_U261 : XNOR2_X2 port map( A => x_vector_28_port, B => 
                           x_vector_27_port, ZN => mult_42_I3_n338);
   mult_42_I3_U260 : XNOR2_X2 port map( A => x_vector_26_port, B => 
                           x_vector_25_port, ZN => mult_42_I3_n327);
   mult_42_I3_U259 : XNOR2_X2 port map( A => x_vector_24_port, B => 
                           x_vector_23_port, ZN => mult_42_I3_n332);
   mult_42_I3_U258 : INV_X1 port map( A => B(21), ZN => mult_42_I3_n312);
   mult_42_I3_U257 : INV_X1 port map( A => B(20), ZN => mult_42_I3_n313);
   mult_42_I3_U256 : INV_X1 port map( A => x_vector_23_port, ZN => 
                           mult_42_I3_n317);
   mult_42_I3_U255 : INV_X1 port map( A => x_vector_20_port, ZN => 
                           mult_42_I3_n320);
   mult_42_I3_U254 : INV_X1 port map( A => x_vector_27_port, ZN => 
                           mult_42_I3_n315);
   mult_42_I3_U253 : INV_X1 port map( A => x_vector_25_port, ZN => 
                           mult_42_I3_n316);
   mult_42_I3_U252 : INV_X1 port map( A => x_vector_29_port, ZN => 
                           mult_42_I3_n314);
   mult_42_I3_U251 : INV_X1 port map( A => mult_42_I3_n367, ZN => 
                           mult_42_I3_n298);
   mult_42_I3_U250 : INV_X1 port map( A => mult_42_I3_n374, ZN => 
                           mult_42_I3_n300);
   mult_42_I3_U249 : INV_X1 port map( A => mult_42_I3_n25, ZN => 
                           mult_42_I3_n301);
   mult_42_I3_U248 : INV_X1 port map( A => mult_42_I3_n35, ZN => 
                           mult_42_I3_n299);
   mult_42_I3_U247 : INV_X1 port map( A => mult_42_I3_n90, ZN => 
                           mult_42_I3_n311);
   mult_42_I3_U246 : INV_X1 port map( A => mult_42_I3_n50, ZN => 
                           mult_42_I3_n297);
   mult_42_I3_U245 : INV_X1 port map( A => mult_42_I3_n349, ZN => 
                           mult_42_I3_n295);
   mult_42_I3_U244 : INV_X1 port map( A => mult_42_I3_n383, ZN => 
                           mult_42_I3_n302);
   mult_42_I3_U243 : INV_X1 port map( A => mult_42_I3_n351, ZN => 
                           mult_42_I3_n318);
   mult_42_I3_U242 : INV_X1 port map( A => mult_42_I3_n352, ZN => 
                           mult_42_I3_n319);
   mult_42_I3_U241 : INV_X1 port map( A => mult_42_I3_n324, ZN => 
                           mult_42_I3_n306);
   mult_42_I3_U240 : INV_X1 port map( A => mult_42_I3_n84, ZN => 
                           mult_42_I3_n308);
   mult_42_I3_U239 : INV_X1 port map( A => mult_42_I3_n87, ZN => 
                           mult_42_I3_n309);
   mult_42_I3_U238 : INV_X1 port map( A => mult_42_I3_n19, ZN => 
                           mult_42_I3_n303);
   mult_42_I3_U237 : INV_X1 port map( A => mult_42_I3_n321, ZN => 
                           mult_42_I3_n310);
   mult_42_I3_U236 : INV_X1 port map( A => mult_42_I3_n1, ZN => N42);
   mult_42_I3_U235 : INV_X1 port map( A => mult_42_I3_n74, ZN => 
                           mult_42_I3_n305);
   mult_42_I3_U234 : INV_X1 port map( A => mult_42_I3_n79, ZN => 
                           mult_42_I3_n307);
   mult_42_I3_U233 : INV_X1 port map( A => mult_42_I3_n60, ZN => 
                           mult_42_I3_n296);
   mult_42_I3_U232 : INV_X1 port map( A => mult_42_I3_n67, ZN => 
                           mult_42_I3_n304);
   mult_42_I3_U56 : HA_X1 port map( A => mult_42_I3_n148, B => mult_42_I3_n157,
                           CO => mult_42_I3_n89, S => mult_42_I3_n90);
   mult_42_I3_U55 : FA_X1 port map( A => mult_42_I3_n156, B => mult_42_I3_n139,
                           CI => mult_42_I3_n147, CO => mult_42_I3_n87, S => 
                           mult_42_I3_n88);
   mult_42_I3_U54 : HA_X1 port map( A => mult_42_I3_n107, B => mult_42_I3_n138,
                           CO => mult_42_I3_n85, S => mult_42_I3_n86);
   mult_42_I3_U53 : FA_X1 port map( A => mult_42_I3_n146, B => mult_42_I3_n155,
                           CI => mult_42_I3_n86, CO => mult_42_I3_n83, S => 
                           mult_42_I3_n84);
   mult_42_I3_U52 : FA_X1 port map( A => mult_42_I3_n154, B => mult_42_I3_n129,
                           CI => mult_42_I3_n145, CO => mult_42_I3_n81, S => 
                           mult_42_I3_n82);
   mult_42_I3_U51 : FA_X1 port map( A => mult_42_I3_n85, B => mult_42_I3_n137, 
                           CI => mult_42_I3_n82, CO => mult_42_I3_n79, S => 
                           mult_42_I3_n80);
   mult_42_I3_U50 : HA_X1 port map( A => mult_42_I3_n106, B => mult_42_I3_n128,
                           CO => mult_42_I3_n77, S => mult_42_I3_n78);
   mult_42_I3_U49 : FA_X1 port map( A => mult_42_I3_n136, B => mult_42_I3_n153,
                           CI => mult_42_I3_n144, CO => mult_42_I3_n75, S => 
                           mult_42_I3_n76);
   mult_42_I3_U48 : FA_X1 port map( A => mult_42_I3_n81, B => mult_42_I3_n78, 
                           CI => mult_42_I3_n76, CO => mult_42_I3_n73, S => 
                           mult_42_I3_n74);
   mult_42_I3_U47 : FA_X1 port map( A => mult_42_I3_n135, B => mult_42_I3_n119,
                           CI => mult_42_I3_n152, CO => mult_42_I3_n71, S => 
                           mult_42_I3_n72);
   mult_42_I3_U46 : FA_X1 port map( A => mult_42_I3_n127, B => mult_42_I3_n143,
                           CI => mult_42_I3_n77, CO => mult_42_I3_n69, S => 
                           mult_42_I3_n70);
   mult_42_I3_U45 : FA_X1 port map( A => mult_42_I3_n72, B => mult_42_I3_n75, 
                           CI => mult_42_I3_n70, CO => mult_42_I3_n67, S => 
                           mult_42_I3_n68);
   mult_42_I3_U44 : HA_X1 port map( A => mult_42_I3_n105, B => mult_42_I3_n118,
                           CO => mult_42_I3_n65, S => mult_42_I3_n66);
   mult_42_I3_U43 : FA_X1 port map( A => mult_42_I3_n126, B => mult_42_I3_n134,
                           CI => mult_42_I3_n142, CO => mult_42_I3_n63, S => 
                           mult_42_I3_n64);
   mult_42_I3_U42 : FA_X1 port map( A => mult_42_I3_n66, B => mult_42_I3_n151, 
                           CI => mult_42_I3_n71, CO => mult_42_I3_n61, S => 
                           mult_42_I3_n62);
   mult_42_I3_U41 : FA_X1 port map( A => mult_42_I3_n64, B => mult_42_I3_n69, 
                           CI => mult_42_I3_n62, CO => mult_42_I3_n59, S => 
                           mult_42_I3_n60);
   mult_42_I3_U38 : FA_X1 port map( A => mult_42_I3_n133, B => mult_42_I3_n117,
                           CI => mult_42_I3_n295, CO => mult_42_I3_n55, S => 
                           mult_42_I3_n56);
   mult_42_I3_U37 : FA_X1 port map( A => mult_42_I3_n58, B => mult_42_I3_n65, 
                           CI => mult_42_I3_n63, CO => mult_42_I3_n53, S => 
                           mult_42_I3_n54);
   mult_42_I3_U36 : FA_X1 port map( A => mult_42_I3_n61, B => mult_42_I3_n56, 
                           CI => mult_42_I3_n54, CO => mult_42_I3_n51, S => 
                           mult_42_I3_n52);
   mult_42_I3_U34 : FA_X1 port map( A => mult_42_I3_n124, B => mult_42_I3_n116,
                           CI => mult_42_I3_n132, CO => mult_42_I3_n47, S => 
                           mult_42_I3_n48);
   mult_42_I3_U33 : FA_X1 port map( A => mult_42_I3_n57, B => mult_42_I3_n50, 
                           CI => mult_42_I3_n55, CO => mult_42_I3_n45, S => 
                           mult_42_I3_n46);
   mult_42_I3_U32 : FA_X1 port map( A => mult_42_I3_n53, B => mult_42_I3_n48, 
                           CI => mult_42_I3_n46, CO => mult_42_I3_n43, S => 
                           mult_42_I3_n44);
   mult_42_I3_U31 : FA_X1 port map( A => mult_42_I3_n123, B => mult_42_I3_n115,
                           CI => mult_42_I3_n140, CO => mult_42_I3_n41, S => 
                           mult_42_I3_n42);
   mult_42_I3_U30 : FA_X1 port map( A => mult_42_I3_n297, B => mult_42_I3_n131,
                           CI => mult_42_I3_n47, CO => mult_42_I3_n39, S => 
                           mult_42_I3_n40);
   mult_42_I3_U29 : FA_X1 port map( A => mult_42_I3_n45, B => mult_42_I3_n42, 
                           CI => mult_42_I3_n40, CO => mult_42_I3_n37, S => 
                           mult_42_I3_n38);
   mult_42_I3_U27 : FA_X1 port map( A => mult_42_I3_n114, B => mult_42_I3_n122,
                           CI => mult_42_I3_n299, CO => mult_42_I3_n33, S => 
                           mult_42_I3_n34);
   mult_42_I3_U26 : FA_X1 port map( A => mult_42_I3_n34, B => mult_42_I3_n41, 
                           CI => mult_42_I3_n39, CO => mult_42_I3_n31, S => 
                           mult_42_I3_n32);
   mult_42_I3_U25 : FA_X1 port map( A => mult_42_I3_n121, B => mult_42_I3_n35, 
                           CI => mult_42_I3_n298, CO => mult_42_I3_n29, S => 
                           mult_42_I3_n30);
   mult_42_I3_U24 : FA_X1 port map( A => mult_42_I3_n33, B => mult_42_I3_n113, 
                           CI => mult_42_I3_n30, CO => mult_42_I3_n27, S => 
                           mult_42_I3_n28);
   mult_42_I3_U22 : FA_X1 port map( A => mult_42_I3_n301, B => mult_42_I3_n112,
                           CI => mult_42_I3_n29, CO => mult_42_I3_n23, S => 
                           mult_42_I3_n24);
   mult_42_I3_U21 : FA_X1 port map( A => mult_42_I3_n111, B => mult_42_I3_n25, 
                           CI => mult_42_I3_n300, CO => mult_42_I3_n21, S => 
                           mult_42_I3_n22);
   mult_42_I3_U10 : FA_X1 port map( A => mult_42_I3_n52, B => mult_42_I3_n59, 
                           CI => mult_42_I3_n10, CO => mult_42_I3_n9, S => N33)
                           ;
   mult_42_I3_U9 : FA_X1 port map( A => mult_42_I3_n44, B => mult_42_I3_n51, CI
                           => mult_42_I3_n9, CO => mult_42_I3_n8, S => N34);
   mult_42_I3_U8 : FA_X1 port map( A => mult_42_I3_n38, B => mult_42_I3_n43, CI
                           => mult_42_I3_n8, CO => mult_42_I3_n7, S => N35);
   mult_42_I3_U7 : FA_X1 port map( A => mult_42_I3_n32, B => mult_42_I3_n37, CI
                           => mult_42_I3_n7, CO => mult_42_I3_n6, S => N36);
   mult_42_I3_U6 : FA_X1 port map( A => mult_42_I3_n28, B => mult_42_I3_n31, CI
                           => mult_42_I3_n6, CO => mult_42_I3_n5, S => N37);
   mult_42_I3_U5 : FA_X1 port map( A => mult_42_I3_n24, B => mult_42_I3_n27, CI
                           => mult_42_I3_n5, CO => mult_42_I3_n4, S => N38);
   mult_42_I3_U4 : FA_X1 port map( A => mult_42_I3_n23, B => mult_42_I3_n22, CI
                           => mult_42_I3_n4, CO => mult_42_I3_n3, S => N39);
   mult_42_I3_U3 : FA_X1 port map( A => mult_42_I3_n21, B => mult_42_I3_n303, 
                           CI => mult_42_I3_n3, CO => mult_42_I3_n2, S => N40);
   mult_42_I3_U2 : FA_X1 port map( A => mult_42_I3_n302, B => mult_42_I3_n19, 
                           CI => mult_42_I3_n2, CO => mult_42_I3_n1, S => N41);
   mult_42_I4_U391 : NAND2_X1 port map( A1 => x_vector_31_port, A2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n341);
   mult_42_I4_U390 : XNOR2_X1 port map( A => B(32), B => x_vector_31_port, ZN 
                           => mult_42_I4_n340);
   mult_42_I4_U389 : OAI22_X1 port map( A1 => B(31), A2 => mult_42_I4_n341, B1 
                           => mult_42_I4_n340, B2 => mult_42_I4_n320, ZN => 
                           mult_42_I4_n402);
   mult_42_I4_U388 : NAND3_X1 port map( A1 => mult_42_I4_n402, A2 => 
                           mult_42_I4_n312, A3 => x_vector_31_port, ZN => 
                           mult_42_I4_n400);
   mult_42_I4_U387 : XNOR2_X1 port map( A => x_vector_32_port, B => 
                           x_vector_31_port, ZN => mult_42_I4_n352);
   mult_42_I4_U386 : NAND2_X1 port map( A1 => mult_42_I4_n319, A2 => 
                           mult_42_I4_n402, ZN => mult_42_I4_n401);
   mult_42_I4_U385 : MUX2_X1 port map( A => mult_42_I4_n400, B => 
                           mult_42_I4_n401, S => B(30), Z => mult_42_I4_n396);
   mult_42_I4_U384 : XOR2_X1 port map( A => x_vector_33_port, B => 
                           x_vector_32_port, Z => mult_42_I4_n399);
   mult_42_I4_U383 : NAND2_X1 port map( A1 => mult_42_I4_n352, A2 => 
                           mult_42_I4_n399, ZN => mult_42_I4_n351);
   mult_42_I4_U382 : NOR3_X1 port map( A1 => mult_42_I4_n352, A2 => B(30), A3 
                           => mult_42_I4_n317, ZN => mult_42_I4_n398);
   mult_42_I4_U381 : AOI21_X1 port map( B1 => x_vector_33_port, B2 => 
                           mult_42_I4_n318, A => mult_42_I4_n398, ZN => 
                           mult_42_I4_n397);
   mult_42_I4_U380 : OAI222_X1 port map( A1 => mult_42_I4_n396, A2 => 
                           mult_42_I4_n311, B1 => mult_42_I4_n397, B2 => 
                           mult_42_I4_n396, C1 => mult_42_I4_n397, C2 => 
                           mult_42_I4_n311, ZN => mult_42_I4_n395);
   mult_42_I4_U379 : AOI222_X1 port map( A1 => mult_42_I4_n395, A2 => 
                           mult_42_I4_n88, B1 => mult_42_I4_n395, B2 => 
                           mult_42_I4_n89, C1 => mult_42_I4_n89, C2 => 
                           mult_42_I4_n88, ZN => mult_42_I4_n394);
   mult_42_I4_U378 : OAI222_X1 port map( A1 => mult_42_I4_n394, A2 => 
                           mult_42_I4_n308, B1 => mult_42_I4_n394, B2 => 
                           mult_42_I4_n309, C1 => mult_42_I4_n309, C2 => 
                           mult_42_I4_n308, ZN => mult_42_I4_n393);
   mult_42_I4_U377 : AOI222_X1 port map( A1 => mult_42_I4_n393, A2 => 
                           mult_42_I4_n80, B1 => mult_42_I4_n393, B2 => 
                           mult_42_I4_n83, C1 => mult_42_I4_n83, C2 => 
                           mult_42_I4_n80, ZN => mult_42_I4_n392);
   mult_42_I4_U376 : OAI222_X1 port map( A1 => mult_42_I4_n392, A2 => 
                           mult_42_I4_n305, B1 => mult_42_I4_n392, B2 => 
                           mult_42_I4_n307, C1 => mult_42_I4_n307, C2 => 
                           mult_42_I4_n305, ZN => mult_42_I4_n391);
   mult_42_I4_U375 : AOI222_X1 port map( A1 => mult_42_I4_n391, A2 => 
                           mult_42_I4_n68, B1 => mult_42_I4_n391, B2 => 
                           mult_42_I4_n73, C1 => mult_42_I4_n73, C2 => 
                           mult_42_I4_n68, ZN => mult_42_I4_n390);
   mult_42_I4_U374 : OAI222_X1 port map( A1 => mult_42_I4_n390, A2 => 
                           mult_42_I4_n296, B1 => mult_42_I4_n390, B2 => 
                           mult_42_I4_n304, C1 => mult_42_I4_n304, C2 => 
                           mult_42_I4_n296, ZN => mult_42_I4_n10);
   mult_42_I4_U373 : XOR2_X1 port map( A => x_vector_39_port, B => 
                           x_vector_38_port, Z => mult_42_I4_n389);
   mult_42_I4_U372 : NAND2_X1 port map( A1 => mult_42_I4_n338, A2 => 
                           mult_42_I4_n389, ZN => mult_42_I4_n337);
   mult_42_I4_U371 : OR3_X1 port map( A1 => mult_42_I4_n338, A2 => B(30), A3 =>
                           mult_42_I4_n314, ZN => mult_42_I4_n388);
   mult_42_I4_U370 : OAI21_X1 port map( B1 => mult_42_I4_n314, B2 => 
                           mult_42_I4_n337, A => mult_42_I4_n388, ZN => 
                           mult_42_I4_n105);
   mult_42_I4_U369 : XOR2_X1 port map( A => x_vector_37_port, B => 
                           x_vector_36_port, Z => mult_42_I4_n387);
   mult_42_I4_U368 : NAND2_X1 port map( A1 => mult_42_I4_n327, A2 => 
                           mult_42_I4_n387, ZN => mult_42_I4_n326);
   mult_42_I4_U367 : OR3_X1 port map( A1 => mult_42_I4_n327, A2 => B(30), A3 =>
                           mult_42_I4_n315, ZN => mult_42_I4_n386);
   mult_42_I4_U366 : OAI21_X1 port map( B1 => mult_42_I4_n315, B2 => 
                           mult_42_I4_n326, A => mult_42_I4_n386, ZN => 
                           mult_42_I4_n106);
   mult_42_I4_U365 : XOR2_X1 port map( A => x_vector_35_port, B => 
                           x_vector_34_port, Z => mult_42_I4_n385);
   mult_42_I4_U364 : NAND2_X1 port map( A1 => mult_42_I4_n332, A2 => 
                           mult_42_I4_n385, ZN => mult_42_I4_n331);
   mult_42_I4_U363 : OR3_X1 port map( A1 => mult_42_I4_n332, A2 => B(30), A3 =>
                           mult_42_I4_n316, ZN => mult_42_I4_n384);
   mult_42_I4_U362 : OAI21_X1 port map( B1 => mult_42_I4_n316, B2 => 
                           mult_42_I4_n331, A => mult_42_I4_n384, ZN => 
                           mult_42_I4_n107);
   mult_42_I4_U361 : XOR2_X1 port map( A => B(39), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n339);
   mult_42_I4_U360 : OAI22_X1 port map( A1 => mult_42_I4_n339, A2 => 
                           mult_42_I4_n338, B1 => mult_42_I4_n337, B2 => 
                           mult_42_I4_n339, ZN => mult_42_I4_n383);
   mult_42_I4_U359 : XOR2_X1 port map( A => B(37), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n382);
   mult_42_I4_U358 : XOR2_X1 port map( A => B(38), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n336);
   mult_42_I4_U357 : OAI22_X1 port map( A1 => mult_42_I4_n382, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n336, ZN => mult_42_I4_n111);
   mult_42_I4_U356 : XOR2_X1 port map( A => B(36), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n381);
   mult_42_I4_U355 : OAI22_X1 port map( A1 => mult_42_I4_n381, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n382, ZN => mult_42_I4_n112);
   mult_42_I4_U354 : XOR2_X1 port map( A => B(35), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n380);
   mult_42_I4_U353 : OAI22_X1 port map( A1 => mult_42_I4_n380, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n381, ZN => mult_42_I4_n113);
   mult_42_I4_U352 : XOR2_X1 port map( A => B(34), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n379);
   mult_42_I4_U351 : OAI22_X1 port map( A1 => mult_42_I4_n379, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n380, ZN => mult_42_I4_n114);
   mult_42_I4_U350 : XOR2_X1 port map( A => B(33), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n378);
   mult_42_I4_U349 : OAI22_X1 port map( A1 => mult_42_I4_n378, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n379, ZN => mult_42_I4_n115);
   mult_42_I4_U348 : XOR2_X1 port map( A => B(32), B => mult_42_I4_n314, Z => 
                           mult_42_I4_n377);
   mult_42_I4_U347 : OAI22_X1 port map( A1 => mult_42_I4_n377, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n378, ZN => mult_42_I4_n116);
   mult_42_I4_U346 : XOR2_X1 port map( A => mult_42_I4_n312, B => 
                           x_vector_39_port, Z => mult_42_I4_n376);
   mult_42_I4_U345 : OAI22_X1 port map( A1 => mult_42_I4_n376, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n377, ZN => mult_42_I4_n117);
   mult_42_I4_U344 : XOR2_X1 port map( A => mult_42_I4_n314, B => B(30), Z => 
                           mult_42_I4_n375);
   mult_42_I4_U343 : OAI22_X1 port map( A1 => mult_42_I4_n375, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n376, ZN => mult_42_I4_n118);
   mult_42_I4_U342 : NOR2_X1 port map( A1 => mult_42_I4_n338, A2 => 
                           mult_42_I4_n313, ZN => mult_42_I4_n119);
   mult_42_I4_U341 : XOR2_X1 port map( A => B(39), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n335);
   mult_42_I4_U340 : OAI22_X1 port map( A1 => mult_42_I4_n335, A2 => 
                           mult_42_I4_n327, B1 => mult_42_I4_n326, B2 => 
                           mult_42_I4_n335, ZN => mult_42_I4_n374);
   mult_42_I4_U339 : XOR2_X1 port map( A => B(37), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n373);
   mult_42_I4_U338 : XOR2_X1 port map( A => B(38), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n334);
   mult_42_I4_U337 : OAI22_X1 port map( A1 => mult_42_I4_n373, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n334, ZN => mult_42_I4_n121);
   mult_42_I4_U336 : XOR2_X1 port map( A => B(36), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n372);
   mult_42_I4_U335 : OAI22_X1 port map( A1 => mult_42_I4_n372, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n373, ZN => mult_42_I4_n122);
   mult_42_I4_U334 : XOR2_X1 port map( A => B(35), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n371);
   mult_42_I4_U333 : OAI22_X1 port map( A1 => mult_42_I4_n371, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n372, ZN => mult_42_I4_n123);
   mult_42_I4_U332 : XOR2_X1 port map( A => B(34), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n328);
   mult_42_I4_U331 : OAI22_X1 port map( A1 => mult_42_I4_n328, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n371, ZN => mult_42_I4_n124);
   mult_42_I4_U330 : XOR2_X1 port map( A => B(32), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n370);
   mult_42_I4_U329 : XOR2_X1 port map( A => B(33), B => mult_42_I4_n315, Z => 
                           mult_42_I4_n325);
   mult_42_I4_U328 : OAI22_X1 port map( A1 => mult_42_I4_n370, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n325, ZN => mult_42_I4_n126);
   mult_42_I4_U327 : XOR2_X1 port map( A => mult_42_I4_n312, B => 
                           x_vector_37_port, Z => mult_42_I4_n369);
   mult_42_I4_U326 : OAI22_X1 port map( A1 => mult_42_I4_n369, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n370, ZN => mult_42_I4_n127);
   mult_42_I4_U325 : XOR2_X1 port map( A => mult_42_I4_n313, B => 
                           x_vector_37_port, Z => mult_42_I4_n368);
   mult_42_I4_U324 : OAI22_X1 port map( A1 => mult_42_I4_n368, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n369, ZN => mult_42_I4_n128);
   mult_42_I4_U323 : NOR2_X1 port map( A1 => mult_42_I4_n327, A2 => 
                           mult_42_I4_n313, ZN => mult_42_I4_n129);
   mult_42_I4_U322 : XOR2_X1 port map( A => B(39), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n333);
   mult_42_I4_U321 : OAI22_X1 port map( A1 => mult_42_I4_n333, A2 => 
                           mult_42_I4_n332, B1 => mult_42_I4_n331, B2 => 
                           mult_42_I4_n333, ZN => mult_42_I4_n367);
   mult_42_I4_U320 : XOR2_X1 port map( A => B(37), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n366);
   mult_42_I4_U319 : XOR2_X1 port map( A => B(38), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n330);
   mult_42_I4_U318 : OAI22_X1 port map( A1 => mult_42_I4_n366, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n330, ZN => mult_42_I4_n131);
   mult_42_I4_U317 : XOR2_X1 port map( A => B(36), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n365);
   mult_42_I4_U316 : OAI22_X1 port map( A1 => mult_42_I4_n365, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n366, ZN => mult_42_I4_n132);
   mult_42_I4_U315 : XOR2_X1 port map( A => B(35), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n364);
   mult_42_I4_U314 : OAI22_X1 port map( A1 => mult_42_I4_n364, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n365, ZN => mult_42_I4_n133);
   mult_42_I4_U313 : XOR2_X1 port map( A => B(34), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n363);
   mult_42_I4_U312 : OAI22_X1 port map( A1 => mult_42_I4_n363, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n364, ZN => mult_42_I4_n134);
   mult_42_I4_U311 : XOR2_X1 port map( A => B(33), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n362);
   mult_42_I4_U310 : OAI22_X1 port map( A1 => mult_42_I4_n362, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n363, ZN => mult_42_I4_n135);
   mult_42_I4_U309 : XOR2_X1 port map( A => B(32), B => mult_42_I4_n316, Z => 
                           mult_42_I4_n361);
   mult_42_I4_U308 : OAI22_X1 port map( A1 => mult_42_I4_n361, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n362, ZN => mult_42_I4_n136);
   mult_42_I4_U307 : XOR2_X1 port map( A => mult_42_I4_n312, B => 
                           x_vector_35_port, Z => mult_42_I4_n360);
   mult_42_I4_U306 : OAI22_X1 port map( A1 => mult_42_I4_n360, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n361, ZN => mult_42_I4_n137);
   mult_42_I4_U305 : XOR2_X1 port map( A => mult_42_I4_n313, B => 
                           x_vector_35_port, Z => mult_42_I4_n359);
   mult_42_I4_U304 : OAI22_X1 port map( A1 => mult_42_I4_n359, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n360, ZN => mult_42_I4_n138);
   mult_42_I4_U303 : NOR2_X1 port map( A1 => mult_42_I4_n332, A2 => 
                           mult_42_I4_n313, ZN => mult_42_I4_n139);
   mult_42_I4_U302 : XOR2_X1 port map( A => B(39), B => x_vector_33_port, Z => 
                           mult_42_I4_n329);
   mult_42_I4_U301 : AOI22_X1 port map( A1 => mult_42_I4_n329, A2 => 
                           mult_42_I4_n319, B1 => mult_42_I4_n318, B2 => 
                           mult_42_I4_n329, ZN => mult_42_I4_n140);
   mult_42_I4_U300 : XOR2_X1 port map( A => B(36), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n358);
   mult_42_I4_U299 : XOR2_X1 port map( A => B(37), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n324);
   mult_42_I4_U298 : OAI22_X1 port map( A1 => mult_42_I4_n358, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n324, ZN => mult_42_I4_n142);
   mult_42_I4_U297 : XOR2_X1 port map( A => B(35), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n357);
   mult_42_I4_U296 : OAI22_X1 port map( A1 => mult_42_I4_n357, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n358, ZN => mult_42_I4_n143);
   mult_42_I4_U295 : XOR2_X1 port map( A => B(34), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n356);
   mult_42_I4_U294 : OAI22_X1 port map( A1 => mult_42_I4_n356, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n357, ZN => mult_42_I4_n144);
   mult_42_I4_U293 : XOR2_X1 port map( A => B(33), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n355);
   mult_42_I4_U292 : OAI22_X1 port map( A1 => mult_42_I4_n355, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n356, ZN => mult_42_I4_n145);
   mult_42_I4_U291 : XOR2_X1 port map( A => B(32), B => mult_42_I4_n317, Z => 
                           mult_42_I4_n354);
   mult_42_I4_U290 : OAI22_X1 port map( A1 => mult_42_I4_n354, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n355, ZN => mult_42_I4_n146);
   mult_42_I4_U289 : XOR2_X1 port map( A => mult_42_I4_n312, B => 
                           x_vector_33_port, Z => mult_42_I4_n353);
   mult_42_I4_U288 : OAI22_X1 port map( A1 => mult_42_I4_n353, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n354, ZN => mult_42_I4_n147);
   mult_42_I4_U287 : XOR2_X1 port map( A => mult_42_I4_n313, B => 
                           x_vector_33_port, Z => mult_42_I4_n350);
   mult_42_I4_U286 : OAI22_X1 port map( A1 => mult_42_I4_n350, A2 => 
                           mult_42_I4_n351, B1 => mult_42_I4_n352, B2 => 
                           mult_42_I4_n353, ZN => mult_42_I4_n148);
   mult_42_I4_U285 : XNOR2_X1 port map( A => B(39), B => x_vector_31_port, ZN 
                           => mult_42_I4_n348);
   mult_42_I4_U284 : OAI22_X1 port map( A1 => mult_42_I4_n320, A2 => 
                           mult_42_I4_n348, B1 => mult_42_I4_n341, B2 => 
                           mult_42_I4_n348, ZN => mult_42_I4_n349);
   mult_42_I4_U283 : XNOR2_X1 port map( A => B(38), B => x_vector_31_port, ZN 
                           => mult_42_I4_n347);
   mult_42_I4_U282 : OAI22_X1 port map( A1 => mult_42_I4_n347, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n348, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n151);
   mult_42_I4_U281 : XNOR2_X1 port map( A => B(37), B => x_vector_31_port, ZN 
                           => mult_42_I4_n346);
   mult_42_I4_U280 : OAI22_X1 port map( A1 => mult_42_I4_n346, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n347, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n152);
   mult_42_I4_U279 : XNOR2_X1 port map( A => B(36), B => x_vector_31_port, ZN 
                           => mult_42_I4_n345);
   mult_42_I4_U278 : OAI22_X1 port map( A1 => mult_42_I4_n345, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n346, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n153);
   mult_42_I4_U277 : XNOR2_X1 port map( A => B(35), B => x_vector_31_port, ZN 
                           => mult_42_I4_n344);
   mult_42_I4_U276 : OAI22_X1 port map( A1 => mult_42_I4_n344, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n345, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n154);
   mult_42_I4_U275 : XNOR2_X1 port map( A => B(34), B => x_vector_31_port, ZN 
                           => mult_42_I4_n343);
   mult_42_I4_U274 : OAI22_X1 port map( A1 => mult_42_I4_n343, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n344, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n155);
   mult_42_I4_U273 : XNOR2_X1 port map( A => B(33), B => x_vector_31_port, ZN 
                           => mult_42_I4_n342);
   mult_42_I4_U272 : OAI22_X1 port map( A1 => mult_42_I4_n342, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n343, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n156);
   mult_42_I4_U271 : OAI22_X1 port map( A1 => mult_42_I4_n340, A2 => 
                           mult_42_I4_n341, B1 => mult_42_I4_n342, B2 => 
                           mult_42_I4_n320, ZN => mult_42_I4_n157);
   mult_42_I4_U270 : OAI22_X1 port map( A1 => mult_42_I4_n336, A2 => 
                           mult_42_I4_n337, B1 => mult_42_I4_n338, B2 => 
                           mult_42_I4_n339, ZN => mult_42_I4_n19);
   mult_42_I4_U269 : OAI22_X1 port map( A1 => mult_42_I4_n334, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n335, ZN => mult_42_I4_n25);
   mult_42_I4_U268 : OAI22_X1 port map( A1 => mult_42_I4_n330, A2 => 
                           mult_42_I4_n331, B1 => mult_42_I4_n332, B2 => 
                           mult_42_I4_n333, ZN => mult_42_I4_n35);
   mult_42_I4_U267 : XOR2_X1 port map( A => B(38), B => x_vector_33_port, Z => 
                           mult_42_I4_n323);
   mult_42_I4_U266 : AOI22_X1 port map( A1 => mult_42_I4_n323, A2 => 
                           mult_42_I4_n318, B1 => mult_42_I4_n319, B2 => 
                           mult_42_I4_n329, ZN => mult_42_I4_n50);
   mult_42_I4_U265 : OAI22_X1 port map( A1 => mult_42_I4_n325, A2 => 
                           mult_42_I4_n326, B1 => mult_42_I4_n327, B2 => 
                           mult_42_I4_n328, ZN => mult_42_I4_n321);
   mult_42_I4_U264 : AOI22_X1 port map( A1 => mult_42_I4_n306, A2 => 
                           mult_42_I4_n318, B1 => mult_42_I4_n319, B2 => 
                           mult_42_I4_n323, ZN => mult_42_I4_n322);
   mult_42_I4_U263 : NAND2_X1 port map( A1 => mult_42_I4_n310, A2 => 
                           mult_42_I4_n322, ZN => mult_42_I4_n57);
   mult_42_I4_U262 : XOR2_X1 port map( A => mult_42_I4_n321, B => 
                           mult_42_I4_n322, Z => mult_42_I4_n58);
   mult_42_I4_U261 : XNOR2_X2 port map( A => x_vector_38_port, B => 
                           x_vector_37_port, ZN => mult_42_I4_n338);
   mult_42_I4_U260 : XNOR2_X2 port map( A => x_vector_36_port, B => 
                           x_vector_35_port, ZN => mult_42_I4_n327);
   mult_42_I4_U259 : XNOR2_X2 port map( A => x_vector_34_port, B => 
                           x_vector_33_port, ZN => mult_42_I4_n332);
   mult_42_I4_U258 : INV_X1 port map( A => B(31), ZN => mult_42_I4_n312);
   mult_42_I4_U257 : INV_X1 port map( A => B(30), ZN => mult_42_I4_n313);
   mult_42_I4_U256 : INV_X1 port map( A => x_vector_33_port, ZN => 
                           mult_42_I4_n317);
   mult_42_I4_U255 : INV_X1 port map( A => x_vector_30_port, ZN => 
                           mult_42_I4_n320);
   mult_42_I4_U254 : INV_X1 port map( A => x_vector_37_port, ZN => 
                           mult_42_I4_n315);
   mult_42_I4_U253 : INV_X1 port map( A => x_vector_35_port, ZN => 
                           mult_42_I4_n316);
   mult_42_I4_U252 : INV_X1 port map( A => x_vector_39_port, ZN => 
                           mult_42_I4_n314);
   mult_42_I4_U251 : INV_X1 port map( A => mult_42_I4_n367, ZN => 
                           mult_42_I4_n298);
   mult_42_I4_U250 : INV_X1 port map( A => mult_42_I4_n374, ZN => 
                           mult_42_I4_n300);
   mult_42_I4_U249 : INV_X1 port map( A => mult_42_I4_n25, ZN => 
                           mult_42_I4_n301);
   mult_42_I4_U248 : INV_X1 port map( A => mult_42_I4_n35, ZN => 
                           mult_42_I4_n299);
   mult_42_I4_U247 : INV_X1 port map( A => mult_42_I4_n90, ZN => 
                           mult_42_I4_n311);
   mult_42_I4_U246 : INV_X1 port map( A => mult_42_I4_n50, ZN => 
                           mult_42_I4_n297);
   mult_42_I4_U245 : INV_X1 port map( A => mult_42_I4_n383, ZN => 
                           mult_42_I4_n302);
   mult_42_I4_U244 : INV_X1 port map( A => mult_42_I4_n349, ZN => 
                           mult_42_I4_n295);
   mult_42_I4_U243 : INV_X1 port map( A => mult_42_I4_n351, ZN => 
                           mult_42_I4_n318);
   mult_42_I4_U242 : INV_X1 port map( A => mult_42_I4_n352, ZN => 
                           mult_42_I4_n319);
   mult_42_I4_U241 : INV_X1 port map( A => mult_42_I4_n324, ZN => 
                           mult_42_I4_n306);
   mult_42_I4_U240 : INV_X1 port map( A => mult_42_I4_n84, ZN => 
                           mult_42_I4_n308);
   mult_42_I4_U239 : INV_X1 port map( A => mult_42_I4_n87, ZN => 
                           mult_42_I4_n309);
   mult_42_I4_U238 : INV_X1 port map( A => mult_42_I4_n19, ZN => 
                           mult_42_I4_n303);
   mult_42_I4_U237 : INV_X1 port map( A => mult_42_I4_n321, ZN => 
                           mult_42_I4_n310);
   mult_42_I4_U236 : INV_X1 port map( A => mult_42_I4_n1, ZN => N62);
   mult_42_I4_U235 : INV_X1 port map( A => mult_42_I4_n74, ZN => 
                           mult_42_I4_n305);
   mult_42_I4_U234 : INV_X1 port map( A => mult_42_I4_n79, ZN => 
                           mult_42_I4_n307);
   mult_42_I4_U233 : INV_X1 port map( A => mult_42_I4_n60, ZN => 
                           mult_42_I4_n296);
   mult_42_I4_U232 : INV_X1 port map( A => mult_42_I4_n67, ZN => 
                           mult_42_I4_n304);
   mult_42_I4_U56 : HA_X1 port map( A => mult_42_I4_n148, B => mult_42_I4_n157,
                           CO => mult_42_I4_n89, S => mult_42_I4_n90);
   mult_42_I4_U55 : FA_X1 port map( A => mult_42_I4_n156, B => mult_42_I4_n139,
                           CI => mult_42_I4_n147, CO => mult_42_I4_n87, S => 
                           mult_42_I4_n88);
   mult_42_I4_U54 : HA_X1 port map( A => mult_42_I4_n107, B => mult_42_I4_n138,
                           CO => mult_42_I4_n85, S => mult_42_I4_n86);
   mult_42_I4_U53 : FA_X1 port map( A => mult_42_I4_n146, B => mult_42_I4_n155,
                           CI => mult_42_I4_n86, CO => mult_42_I4_n83, S => 
                           mult_42_I4_n84);
   mult_42_I4_U52 : FA_X1 port map( A => mult_42_I4_n154, B => mult_42_I4_n129,
                           CI => mult_42_I4_n145, CO => mult_42_I4_n81, S => 
                           mult_42_I4_n82);
   mult_42_I4_U51 : FA_X1 port map( A => mult_42_I4_n85, B => mult_42_I4_n137, 
                           CI => mult_42_I4_n82, CO => mult_42_I4_n79, S => 
                           mult_42_I4_n80);
   mult_42_I4_U50 : HA_X1 port map( A => mult_42_I4_n106, B => mult_42_I4_n128,
                           CO => mult_42_I4_n77, S => mult_42_I4_n78);
   mult_42_I4_U49 : FA_X1 port map( A => mult_42_I4_n136, B => mult_42_I4_n153,
                           CI => mult_42_I4_n144, CO => mult_42_I4_n75, S => 
                           mult_42_I4_n76);
   mult_42_I4_U48 : FA_X1 port map( A => mult_42_I4_n81, B => mult_42_I4_n78, 
                           CI => mult_42_I4_n76, CO => mult_42_I4_n73, S => 
                           mult_42_I4_n74);
   mult_42_I4_U47 : FA_X1 port map( A => mult_42_I4_n135, B => mult_42_I4_n119,
                           CI => mult_42_I4_n152, CO => mult_42_I4_n71, S => 
                           mult_42_I4_n72);
   mult_42_I4_U46 : FA_X1 port map( A => mult_42_I4_n127, B => mult_42_I4_n143,
                           CI => mult_42_I4_n77, CO => mult_42_I4_n69, S => 
                           mult_42_I4_n70);
   mult_42_I4_U45 : FA_X1 port map( A => mult_42_I4_n72, B => mult_42_I4_n75, 
                           CI => mult_42_I4_n70, CO => mult_42_I4_n67, S => 
                           mult_42_I4_n68);
   mult_42_I4_U44 : HA_X1 port map( A => mult_42_I4_n105, B => mult_42_I4_n118,
                           CO => mult_42_I4_n65, S => mult_42_I4_n66);
   mult_42_I4_U43 : FA_X1 port map( A => mult_42_I4_n126, B => mult_42_I4_n134,
                           CI => mult_42_I4_n142, CO => mult_42_I4_n63, S => 
                           mult_42_I4_n64);
   mult_42_I4_U42 : FA_X1 port map( A => mult_42_I4_n66, B => mult_42_I4_n151, 
                           CI => mult_42_I4_n71, CO => mult_42_I4_n61, S => 
                           mult_42_I4_n62);
   mult_42_I4_U41 : FA_X1 port map( A => mult_42_I4_n64, B => mult_42_I4_n69, 
                           CI => mult_42_I4_n62, CO => mult_42_I4_n59, S => 
                           mult_42_I4_n60);
   mult_42_I4_U38 : FA_X1 port map( A => mult_42_I4_n133, B => mult_42_I4_n117,
                           CI => mult_42_I4_n295, CO => mult_42_I4_n55, S => 
                           mult_42_I4_n56);
   mult_42_I4_U37 : FA_X1 port map( A => mult_42_I4_n58, B => mult_42_I4_n65, 
                           CI => mult_42_I4_n63, CO => mult_42_I4_n53, S => 
                           mult_42_I4_n54);
   mult_42_I4_U36 : FA_X1 port map( A => mult_42_I4_n61, B => mult_42_I4_n56, 
                           CI => mult_42_I4_n54, CO => mult_42_I4_n51, S => 
                           mult_42_I4_n52);
   mult_42_I4_U34 : FA_X1 port map( A => mult_42_I4_n124, B => mult_42_I4_n116,
                           CI => mult_42_I4_n132, CO => mult_42_I4_n47, S => 
                           mult_42_I4_n48);
   mult_42_I4_U33 : FA_X1 port map( A => mult_42_I4_n57, B => mult_42_I4_n50, 
                           CI => mult_42_I4_n55, CO => mult_42_I4_n45, S => 
                           mult_42_I4_n46);
   mult_42_I4_U32 : FA_X1 port map( A => mult_42_I4_n53, B => mult_42_I4_n48, 
                           CI => mult_42_I4_n46, CO => mult_42_I4_n43, S => 
                           mult_42_I4_n44);
   mult_42_I4_U31 : FA_X1 port map( A => mult_42_I4_n123, B => mult_42_I4_n115,
                           CI => mult_42_I4_n140, CO => mult_42_I4_n41, S => 
                           mult_42_I4_n42);
   mult_42_I4_U30 : FA_X1 port map( A => mult_42_I4_n297, B => mult_42_I4_n131,
                           CI => mult_42_I4_n47, CO => mult_42_I4_n39, S => 
                           mult_42_I4_n40);
   mult_42_I4_U29 : FA_X1 port map( A => mult_42_I4_n45, B => mult_42_I4_n42, 
                           CI => mult_42_I4_n40, CO => mult_42_I4_n37, S => 
                           mult_42_I4_n38);
   mult_42_I4_U27 : FA_X1 port map( A => mult_42_I4_n114, B => mult_42_I4_n122,
                           CI => mult_42_I4_n299, CO => mult_42_I4_n33, S => 
                           mult_42_I4_n34);
   mult_42_I4_U26 : FA_X1 port map( A => mult_42_I4_n34, B => mult_42_I4_n41, 
                           CI => mult_42_I4_n39, CO => mult_42_I4_n31, S => 
                           mult_42_I4_n32);
   mult_42_I4_U25 : FA_X1 port map( A => mult_42_I4_n121, B => mult_42_I4_n35, 
                           CI => mult_42_I4_n298, CO => mult_42_I4_n29, S => 
                           mult_42_I4_n30);
   mult_42_I4_U24 : FA_X1 port map( A => mult_42_I4_n33, B => mult_42_I4_n113, 
                           CI => mult_42_I4_n30, CO => mult_42_I4_n27, S => 
                           mult_42_I4_n28);
   mult_42_I4_U22 : FA_X1 port map( A => mult_42_I4_n301, B => mult_42_I4_n112,
                           CI => mult_42_I4_n29, CO => mult_42_I4_n23, S => 
                           mult_42_I4_n24);
   mult_42_I4_U21 : FA_X1 port map( A => mult_42_I4_n111, B => mult_42_I4_n25, 
                           CI => mult_42_I4_n300, CO => mult_42_I4_n21, S => 
                           mult_42_I4_n22);
   mult_42_I4_U10 : FA_X1 port map( A => mult_42_I4_n52, B => mult_42_I4_n59, 
                           CI => mult_42_I4_n10, CO => mult_42_I4_n9, S => N53)
                           ;
   mult_42_I4_U9 : FA_X1 port map( A => mult_42_I4_n44, B => mult_42_I4_n51, CI
                           => mult_42_I4_n9, CO => mult_42_I4_n8, S => N54);
   mult_42_I4_U8 : FA_X1 port map( A => mult_42_I4_n38, B => mult_42_I4_n43, CI
                           => mult_42_I4_n8, CO => mult_42_I4_n7, S => N55);
   mult_42_I4_U7 : FA_X1 port map( A => mult_42_I4_n32, B => mult_42_I4_n37, CI
                           => mult_42_I4_n7, CO => mult_42_I4_n6, S => N56);
   mult_42_I4_U6 : FA_X1 port map( A => mult_42_I4_n28, B => mult_42_I4_n31, CI
                           => mult_42_I4_n6, CO => mult_42_I4_n5, S => N57);
   mult_42_I4_U5 : FA_X1 port map( A => mult_42_I4_n24, B => mult_42_I4_n27, CI
                           => mult_42_I4_n5, CO => mult_42_I4_n4, S => N58);
   mult_42_I4_U4 : FA_X1 port map( A => mult_42_I4_n23, B => mult_42_I4_n22, CI
                           => mult_42_I4_n4, CO => mult_42_I4_n3, S => N59);
   mult_42_I4_U3 : FA_X1 port map( A => mult_42_I4_n21, B => mult_42_I4_n303, 
                           CI => mult_42_I4_n3, CO => mult_42_I4_n2, S => N60);
   mult_42_I4_U2 : FA_X1 port map( A => mult_42_I4_n302, B => mult_42_I4_n19, 
                           CI => mult_42_I4_n2, CO => mult_42_I4_n1, S => N61);
   mult_42_I5_U391 : NAND2_X1 port map( A1 => x_vector_41_port, A2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n341);
   mult_42_I5_U390 : XNOR2_X1 port map( A => B(42), B => x_vector_41_port, ZN 
                           => mult_42_I5_n340);
   mult_42_I5_U389 : OAI22_X1 port map( A1 => B(41), A2 => mult_42_I5_n341, B1 
                           => mult_42_I5_n340, B2 => mult_42_I5_n320, ZN => 
                           mult_42_I5_n402);
   mult_42_I5_U388 : NAND3_X1 port map( A1 => mult_42_I5_n402, A2 => 
                           mult_42_I5_n312, A3 => x_vector_41_port, ZN => 
                           mult_42_I5_n400);
   mult_42_I5_U387 : XNOR2_X1 port map( A => x_vector_42_port, B => 
                           x_vector_41_port, ZN => mult_42_I5_n352);
   mult_42_I5_U386 : NAND2_X1 port map( A1 => mult_42_I5_n319, A2 => 
                           mult_42_I5_n402, ZN => mult_42_I5_n401);
   mult_42_I5_U385 : MUX2_X1 port map( A => mult_42_I5_n400, B => 
                           mult_42_I5_n401, S => B(40), Z => mult_42_I5_n396);
   mult_42_I5_U384 : XOR2_X1 port map( A => x_vector_43_port, B => 
                           x_vector_42_port, Z => mult_42_I5_n399);
   mult_42_I5_U383 : NAND2_X1 port map( A1 => mult_42_I5_n352, A2 => 
                           mult_42_I5_n399, ZN => mult_42_I5_n351);
   mult_42_I5_U382 : NOR3_X1 port map( A1 => mult_42_I5_n352, A2 => B(40), A3 
                           => mult_42_I5_n317, ZN => mult_42_I5_n398);
   mult_42_I5_U381 : AOI21_X1 port map( B1 => x_vector_43_port, B2 => 
                           mult_42_I5_n318, A => mult_42_I5_n398, ZN => 
                           mult_42_I5_n397);
   mult_42_I5_U380 : OAI222_X1 port map( A1 => mult_42_I5_n396, A2 => 
                           mult_42_I5_n311, B1 => mult_42_I5_n397, B2 => 
                           mult_42_I5_n396, C1 => mult_42_I5_n397, C2 => 
                           mult_42_I5_n311, ZN => mult_42_I5_n395);
   mult_42_I5_U379 : AOI222_X1 port map( A1 => mult_42_I5_n395, A2 => 
                           mult_42_I5_n88, B1 => mult_42_I5_n395, B2 => 
                           mult_42_I5_n89, C1 => mult_42_I5_n89, C2 => 
                           mult_42_I5_n88, ZN => mult_42_I5_n394);
   mult_42_I5_U378 : OAI222_X1 port map( A1 => mult_42_I5_n394, A2 => 
                           mult_42_I5_n308, B1 => mult_42_I5_n394, B2 => 
                           mult_42_I5_n309, C1 => mult_42_I5_n309, C2 => 
                           mult_42_I5_n308, ZN => mult_42_I5_n393);
   mult_42_I5_U377 : AOI222_X1 port map( A1 => mult_42_I5_n393, A2 => 
                           mult_42_I5_n80, B1 => mult_42_I5_n393, B2 => 
                           mult_42_I5_n83, C1 => mult_42_I5_n83, C2 => 
                           mult_42_I5_n80, ZN => mult_42_I5_n392);
   mult_42_I5_U376 : OAI222_X1 port map( A1 => mult_42_I5_n392, A2 => 
                           mult_42_I5_n305, B1 => mult_42_I5_n392, B2 => 
                           mult_42_I5_n307, C1 => mult_42_I5_n307, C2 => 
                           mult_42_I5_n305, ZN => mult_42_I5_n391);
   mult_42_I5_U375 : AOI222_X1 port map( A1 => mult_42_I5_n391, A2 => 
                           mult_42_I5_n68, B1 => mult_42_I5_n391, B2 => 
                           mult_42_I5_n73, C1 => mult_42_I5_n73, C2 => 
                           mult_42_I5_n68, ZN => mult_42_I5_n390);
   mult_42_I5_U374 : OAI222_X1 port map( A1 => mult_42_I5_n390, A2 => 
                           mult_42_I5_n296, B1 => mult_42_I5_n390, B2 => 
                           mult_42_I5_n304, C1 => mult_42_I5_n304, C2 => 
                           mult_42_I5_n296, ZN => mult_42_I5_n10);
   mult_42_I5_U373 : XOR2_X1 port map( A => x_vector_49_port, B => 
                           x_vector_48_port, Z => mult_42_I5_n389);
   mult_42_I5_U372 : NAND2_X1 port map( A1 => mult_42_I5_n338, A2 => 
                           mult_42_I5_n389, ZN => mult_42_I5_n337);
   mult_42_I5_U371 : OR3_X1 port map( A1 => mult_42_I5_n338, A2 => B(40), A3 =>
                           mult_42_I5_n314, ZN => mult_42_I5_n388);
   mult_42_I5_U370 : OAI21_X1 port map( B1 => mult_42_I5_n314, B2 => 
                           mult_42_I5_n337, A => mult_42_I5_n388, ZN => 
                           mult_42_I5_n105);
   mult_42_I5_U369 : XOR2_X1 port map( A => x_vector_47_port, B => 
                           x_vector_46_port, Z => mult_42_I5_n387);
   mult_42_I5_U368 : NAND2_X1 port map( A1 => mult_42_I5_n327, A2 => 
                           mult_42_I5_n387, ZN => mult_42_I5_n326);
   mult_42_I5_U367 : OR3_X1 port map( A1 => mult_42_I5_n327, A2 => B(40), A3 =>
                           mult_42_I5_n315, ZN => mult_42_I5_n386);
   mult_42_I5_U366 : OAI21_X1 port map( B1 => mult_42_I5_n315, B2 => 
                           mult_42_I5_n326, A => mult_42_I5_n386, ZN => 
                           mult_42_I5_n106);
   mult_42_I5_U365 : XOR2_X1 port map( A => x_vector_45_port, B => 
                           x_vector_44_port, Z => mult_42_I5_n385);
   mult_42_I5_U364 : NAND2_X1 port map( A1 => mult_42_I5_n332, A2 => 
                           mult_42_I5_n385, ZN => mult_42_I5_n331);
   mult_42_I5_U363 : OR3_X1 port map( A1 => mult_42_I5_n332, A2 => B(40), A3 =>
                           mult_42_I5_n316, ZN => mult_42_I5_n384);
   mult_42_I5_U362 : OAI21_X1 port map( B1 => mult_42_I5_n316, B2 => 
                           mult_42_I5_n331, A => mult_42_I5_n384, ZN => 
                           mult_42_I5_n107);
   mult_42_I5_U361 : XOR2_X1 port map( A => B(49), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n339);
   mult_42_I5_U360 : OAI22_X1 port map( A1 => mult_42_I5_n339, A2 => 
                           mult_42_I5_n338, B1 => mult_42_I5_n337, B2 => 
                           mult_42_I5_n339, ZN => mult_42_I5_n383);
   mult_42_I5_U359 : XOR2_X1 port map( A => B(47), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n382);
   mult_42_I5_U358 : XOR2_X1 port map( A => B(48), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n336);
   mult_42_I5_U357 : OAI22_X1 port map( A1 => mult_42_I5_n382, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n336, ZN => mult_42_I5_n111);
   mult_42_I5_U356 : XOR2_X1 port map( A => B(46), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n381);
   mult_42_I5_U355 : OAI22_X1 port map( A1 => mult_42_I5_n381, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n382, ZN => mult_42_I5_n112);
   mult_42_I5_U354 : XOR2_X1 port map( A => B(45), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n380);
   mult_42_I5_U353 : OAI22_X1 port map( A1 => mult_42_I5_n380, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n381, ZN => mult_42_I5_n113);
   mult_42_I5_U352 : XOR2_X1 port map( A => B(44), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n379);
   mult_42_I5_U351 : OAI22_X1 port map( A1 => mult_42_I5_n379, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n380, ZN => mult_42_I5_n114);
   mult_42_I5_U350 : XOR2_X1 port map( A => B(43), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n378);
   mult_42_I5_U349 : OAI22_X1 port map( A1 => mult_42_I5_n378, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n379, ZN => mult_42_I5_n115);
   mult_42_I5_U348 : XOR2_X1 port map( A => B(42), B => mult_42_I5_n314, Z => 
                           mult_42_I5_n377);
   mult_42_I5_U347 : OAI22_X1 port map( A1 => mult_42_I5_n377, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n378, ZN => mult_42_I5_n116);
   mult_42_I5_U346 : XOR2_X1 port map( A => mult_42_I5_n312, B => 
                           x_vector_49_port, Z => mult_42_I5_n376);
   mult_42_I5_U345 : OAI22_X1 port map( A1 => mult_42_I5_n376, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n377, ZN => mult_42_I5_n117);
   mult_42_I5_U344 : XOR2_X1 port map( A => mult_42_I5_n314, B => B(40), Z => 
                           mult_42_I5_n375);
   mult_42_I5_U343 : OAI22_X1 port map( A1 => mult_42_I5_n375, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n376, ZN => mult_42_I5_n118);
   mult_42_I5_U342 : NOR2_X1 port map( A1 => mult_42_I5_n338, A2 => 
                           mult_42_I5_n313, ZN => mult_42_I5_n119);
   mult_42_I5_U341 : XOR2_X1 port map( A => B(49), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n335);
   mult_42_I5_U340 : OAI22_X1 port map( A1 => mult_42_I5_n335, A2 => 
                           mult_42_I5_n327, B1 => mult_42_I5_n326, B2 => 
                           mult_42_I5_n335, ZN => mult_42_I5_n374);
   mult_42_I5_U339 : XOR2_X1 port map( A => B(47), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n373);
   mult_42_I5_U338 : XOR2_X1 port map( A => B(48), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n334);
   mult_42_I5_U337 : OAI22_X1 port map( A1 => mult_42_I5_n373, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n334, ZN => mult_42_I5_n121);
   mult_42_I5_U336 : XOR2_X1 port map( A => B(46), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n372);
   mult_42_I5_U335 : OAI22_X1 port map( A1 => mult_42_I5_n372, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n373, ZN => mult_42_I5_n122);
   mult_42_I5_U334 : XOR2_X1 port map( A => B(45), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n371);
   mult_42_I5_U333 : OAI22_X1 port map( A1 => mult_42_I5_n371, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n372, ZN => mult_42_I5_n123);
   mult_42_I5_U332 : XOR2_X1 port map( A => B(44), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n328);
   mult_42_I5_U331 : OAI22_X1 port map( A1 => mult_42_I5_n328, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n371, ZN => mult_42_I5_n124);
   mult_42_I5_U330 : XOR2_X1 port map( A => B(42), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n370);
   mult_42_I5_U329 : XOR2_X1 port map( A => B(43), B => mult_42_I5_n315, Z => 
                           mult_42_I5_n325);
   mult_42_I5_U328 : OAI22_X1 port map( A1 => mult_42_I5_n370, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n325, ZN => mult_42_I5_n126);
   mult_42_I5_U327 : XOR2_X1 port map( A => mult_42_I5_n312, B => 
                           x_vector_47_port, Z => mult_42_I5_n369);
   mult_42_I5_U326 : OAI22_X1 port map( A1 => mult_42_I5_n369, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n370, ZN => mult_42_I5_n127);
   mult_42_I5_U325 : XOR2_X1 port map( A => mult_42_I5_n313, B => 
                           x_vector_47_port, Z => mult_42_I5_n368);
   mult_42_I5_U324 : OAI22_X1 port map( A1 => mult_42_I5_n368, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n369, ZN => mult_42_I5_n128);
   mult_42_I5_U323 : NOR2_X1 port map( A1 => mult_42_I5_n327, A2 => 
                           mult_42_I5_n313, ZN => mult_42_I5_n129);
   mult_42_I5_U322 : XOR2_X1 port map( A => B(49), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n333);
   mult_42_I5_U321 : OAI22_X1 port map( A1 => mult_42_I5_n333, A2 => 
                           mult_42_I5_n332, B1 => mult_42_I5_n331, B2 => 
                           mult_42_I5_n333, ZN => mult_42_I5_n367);
   mult_42_I5_U320 : XOR2_X1 port map( A => B(47), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n366);
   mult_42_I5_U319 : XOR2_X1 port map( A => B(48), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n330);
   mult_42_I5_U318 : OAI22_X1 port map( A1 => mult_42_I5_n366, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n330, ZN => mult_42_I5_n131);
   mult_42_I5_U317 : XOR2_X1 port map( A => B(46), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n365);
   mult_42_I5_U316 : OAI22_X1 port map( A1 => mult_42_I5_n365, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n366, ZN => mult_42_I5_n132);
   mult_42_I5_U315 : XOR2_X1 port map( A => B(45), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n364);
   mult_42_I5_U314 : OAI22_X1 port map( A1 => mult_42_I5_n364, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n365, ZN => mult_42_I5_n133);
   mult_42_I5_U313 : XOR2_X1 port map( A => B(44), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n363);
   mult_42_I5_U312 : OAI22_X1 port map( A1 => mult_42_I5_n363, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n364, ZN => mult_42_I5_n134);
   mult_42_I5_U311 : XOR2_X1 port map( A => B(43), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n362);
   mult_42_I5_U310 : OAI22_X1 port map( A1 => mult_42_I5_n362, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n363, ZN => mult_42_I5_n135);
   mult_42_I5_U309 : XOR2_X1 port map( A => B(42), B => mult_42_I5_n316, Z => 
                           mult_42_I5_n361);
   mult_42_I5_U308 : OAI22_X1 port map( A1 => mult_42_I5_n361, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n362, ZN => mult_42_I5_n136);
   mult_42_I5_U307 : XOR2_X1 port map( A => mult_42_I5_n312, B => 
                           x_vector_45_port, Z => mult_42_I5_n360);
   mult_42_I5_U306 : OAI22_X1 port map( A1 => mult_42_I5_n360, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n361, ZN => mult_42_I5_n137);
   mult_42_I5_U305 : XOR2_X1 port map( A => mult_42_I5_n313, B => 
                           x_vector_45_port, Z => mult_42_I5_n359);
   mult_42_I5_U304 : OAI22_X1 port map( A1 => mult_42_I5_n359, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n360, ZN => mult_42_I5_n138);
   mult_42_I5_U303 : NOR2_X1 port map( A1 => mult_42_I5_n332, A2 => 
                           mult_42_I5_n313, ZN => mult_42_I5_n139);
   mult_42_I5_U302 : XOR2_X1 port map( A => B(49), B => x_vector_43_port, Z => 
                           mult_42_I5_n329);
   mult_42_I5_U301 : AOI22_X1 port map( A1 => mult_42_I5_n329, A2 => 
                           mult_42_I5_n319, B1 => mult_42_I5_n318, B2 => 
                           mult_42_I5_n329, ZN => mult_42_I5_n140);
   mult_42_I5_U300 : XOR2_X1 port map( A => B(46), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n358);
   mult_42_I5_U299 : XOR2_X1 port map( A => B(47), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n324);
   mult_42_I5_U298 : OAI22_X1 port map( A1 => mult_42_I5_n358, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n324, ZN => mult_42_I5_n142);
   mult_42_I5_U297 : XOR2_X1 port map( A => B(45), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n357);
   mult_42_I5_U296 : OAI22_X1 port map( A1 => mult_42_I5_n357, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n358, ZN => mult_42_I5_n143);
   mult_42_I5_U295 : XOR2_X1 port map( A => B(44), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n356);
   mult_42_I5_U294 : OAI22_X1 port map( A1 => mult_42_I5_n356, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n357, ZN => mult_42_I5_n144);
   mult_42_I5_U293 : XOR2_X1 port map( A => B(43), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n355);
   mult_42_I5_U292 : OAI22_X1 port map( A1 => mult_42_I5_n355, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n356, ZN => mult_42_I5_n145);
   mult_42_I5_U291 : XOR2_X1 port map( A => B(42), B => mult_42_I5_n317, Z => 
                           mult_42_I5_n354);
   mult_42_I5_U290 : OAI22_X1 port map( A1 => mult_42_I5_n354, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n355, ZN => mult_42_I5_n146);
   mult_42_I5_U289 : XOR2_X1 port map( A => mult_42_I5_n312, B => 
                           x_vector_43_port, Z => mult_42_I5_n353);
   mult_42_I5_U288 : OAI22_X1 port map( A1 => mult_42_I5_n353, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n354, ZN => mult_42_I5_n147);
   mult_42_I5_U287 : XOR2_X1 port map( A => mult_42_I5_n313, B => 
                           x_vector_43_port, Z => mult_42_I5_n350);
   mult_42_I5_U286 : OAI22_X1 port map( A1 => mult_42_I5_n350, A2 => 
                           mult_42_I5_n351, B1 => mult_42_I5_n352, B2 => 
                           mult_42_I5_n353, ZN => mult_42_I5_n148);
   mult_42_I5_U285 : XNOR2_X1 port map( A => B(49), B => x_vector_41_port, ZN 
                           => mult_42_I5_n348);
   mult_42_I5_U284 : OAI22_X1 port map( A1 => mult_42_I5_n320, A2 => 
                           mult_42_I5_n348, B1 => mult_42_I5_n341, B2 => 
                           mult_42_I5_n348, ZN => mult_42_I5_n349);
   mult_42_I5_U283 : XNOR2_X1 port map( A => B(48), B => x_vector_41_port, ZN 
                           => mult_42_I5_n347);
   mult_42_I5_U282 : OAI22_X1 port map( A1 => mult_42_I5_n347, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n348, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n151);
   mult_42_I5_U281 : XNOR2_X1 port map( A => B(47), B => x_vector_41_port, ZN 
                           => mult_42_I5_n346);
   mult_42_I5_U280 : OAI22_X1 port map( A1 => mult_42_I5_n346, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n347, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n152);
   mult_42_I5_U279 : XNOR2_X1 port map( A => B(46), B => x_vector_41_port, ZN 
                           => mult_42_I5_n345);
   mult_42_I5_U278 : OAI22_X1 port map( A1 => mult_42_I5_n345, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n346, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n153);
   mult_42_I5_U277 : XNOR2_X1 port map( A => B(45), B => x_vector_41_port, ZN 
                           => mult_42_I5_n344);
   mult_42_I5_U276 : OAI22_X1 port map( A1 => mult_42_I5_n344, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n345, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n154);
   mult_42_I5_U275 : XNOR2_X1 port map( A => B(44), B => x_vector_41_port, ZN 
                           => mult_42_I5_n343);
   mult_42_I5_U274 : OAI22_X1 port map( A1 => mult_42_I5_n343, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n344, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n155);
   mult_42_I5_U273 : XNOR2_X1 port map( A => B(43), B => x_vector_41_port, ZN 
                           => mult_42_I5_n342);
   mult_42_I5_U272 : OAI22_X1 port map( A1 => mult_42_I5_n342, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n343, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n156);
   mult_42_I5_U271 : OAI22_X1 port map( A1 => mult_42_I5_n340, A2 => 
                           mult_42_I5_n341, B1 => mult_42_I5_n342, B2 => 
                           mult_42_I5_n320, ZN => mult_42_I5_n157);
   mult_42_I5_U270 : OAI22_X1 port map( A1 => mult_42_I5_n336, A2 => 
                           mult_42_I5_n337, B1 => mult_42_I5_n338, B2 => 
                           mult_42_I5_n339, ZN => mult_42_I5_n19);
   mult_42_I5_U269 : OAI22_X1 port map( A1 => mult_42_I5_n334, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n335, ZN => mult_42_I5_n25);
   mult_42_I5_U268 : OAI22_X1 port map( A1 => mult_42_I5_n330, A2 => 
                           mult_42_I5_n331, B1 => mult_42_I5_n332, B2 => 
                           mult_42_I5_n333, ZN => mult_42_I5_n35);
   mult_42_I5_U267 : XOR2_X1 port map( A => B(48), B => x_vector_43_port, Z => 
                           mult_42_I5_n323);
   mult_42_I5_U266 : AOI22_X1 port map( A1 => mult_42_I5_n323, A2 => 
                           mult_42_I5_n318, B1 => mult_42_I5_n319, B2 => 
                           mult_42_I5_n329, ZN => mult_42_I5_n50);
   mult_42_I5_U265 : OAI22_X1 port map( A1 => mult_42_I5_n325, A2 => 
                           mult_42_I5_n326, B1 => mult_42_I5_n327, B2 => 
                           mult_42_I5_n328, ZN => mult_42_I5_n321);
   mult_42_I5_U264 : AOI22_X1 port map( A1 => mult_42_I5_n306, A2 => 
                           mult_42_I5_n318, B1 => mult_42_I5_n319, B2 => 
                           mult_42_I5_n323, ZN => mult_42_I5_n322);
   mult_42_I5_U263 : NAND2_X1 port map( A1 => mult_42_I5_n310, A2 => 
                           mult_42_I5_n322, ZN => mult_42_I5_n57);
   mult_42_I5_U262 : XOR2_X1 port map( A => mult_42_I5_n321, B => 
                           mult_42_I5_n322, Z => mult_42_I5_n58);
   mult_42_I5_U261 : XNOR2_X2 port map( A => x_vector_48_port, B => 
                           x_vector_47_port, ZN => mult_42_I5_n338);
   mult_42_I5_U260 : XNOR2_X2 port map( A => x_vector_46_port, B => 
                           x_vector_45_port, ZN => mult_42_I5_n327);
   mult_42_I5_U259 : XNOR2_X2 port map( A => x_vector_44_port, B => 
                           x_vector_43_port, ZN => mult_42_I5_n332);
   mult_42_I5_U258 : INV_X1 port map( A => B(41), ZN => mult_42_I5_n312);
   mult_42_I5_U257 : INV_X1 port map( A => B(40), ZN => mult_42_I5_n313);
   mult_42_I5_U256 : INV_X1 port map( A => x_vector_43_port, ZN => 
                           mult_42_I5_n317);
   mult_42_I5_U255 : INV_X1 port map( A => x_vector_40_port, ZN => 
                           mult_42_I5_n320);
   mult_42_I5_U254 : INV_X1 port map( A => x_vector_47_port, ZN => 
                           mult_42_I5_n315);
   mult_42_I5_U253 : INV_X1 port map( A => x_vector_45_port, ZN => 
                           mult_42_I5_n316);
   mult_42_I5_U252 : INV_X1 port map( A => x_vector_49_port, ZN => 
                           mult_42_I5_n314);
   mult_42_I5_U251 : INV_X1 port map( A => mult_42_I5_n374, ZN => 
                           mult_42_I5_n300);
   mult_42_I5_U250 : INV_X1 port map( A => mult_42_I5_n25, ZN => 
                           mult_42_I5_n301);
   mult_42_I5_U249 : INV_X1 port map( A => mult_42_I5_n90, ZN => 
                           mult_42_I5_n311);
   mult_42_I5_U248 : INV_X1 port map( A => mult_42_I5_n50, ZN => 
                           mult_42_I5_n297);
   mult_42_I5_U247 : INV_X1 port map( A => mult_42_I5_n367, ZN => 
                           mult_42_I5_n298);
   mult_42_I5_U246 : INV_X1 port map( A => mult_42_I5_n383, ZN => 
                           mult_42_I5_n302);
   mult_42_I5_U245 : INV_X1 port map( A => mult_42_I5_n349, ZN => 
                           mult_42_I5_n295);
   mult_42_I5_U244 : INV_X1 port map( A => mult_42_I5_n35, ZN => 
                           mult_42_I5_n299);
   mult_42_I5_U243 : INV_X1 port map( A => mult_42_I5_n351, ZN => 
                           mult_42_I5_n318);
   mult_42_I5_U242 : INV_X1 port map( A => mult_42_I5_n352, ZN => 
                           mult_42_I5_n319);
   mult_42_I5_U241 : INV_X1 port map( A => mult_42_I5_n324, ZN => 
                           mult_42_I5_n306);
   mult_42_I5_U240 : INV_X1 port map( A => mult_42_I5_n84, ZN => 
                           mult_42_I5_n308);
   mult_42_I5_U239 : INV_X1 port map( A => mult_42_I5_n87, ZN => 
                           mult_42_I5_n309);
   mult_42_I5_U238 : INV_X1 port map( A => mult_42_I5_n19, ZN => 
                           mult_42_I5_n303);
   mult_42_I5_U237 : INV_X1 port map( A => mult_42_I5_n321, ZN => 
                           mult_42_I5_n310);
   mult_42_I5_U236 : INV_X1 port map( A => mult_42_I5_n1, ZN => N82);
   mult_42_I5_U235 : INV_X1 port map( A => mult_42_I5_n74, ZN => 
                           mult_42_I5_n305);
   mult_42_I5_U234 : INV_X1 port map( A => mult_42_I5_n79, ZN => 
                           mult_42_I5_n307);
   mult_42_I5_U233 : INV_X1 port map( A => mult_42_I5_n60, ZN => 
                           mult_42_I5_n296);
   mult_42_I5_U232 : INV_X1 port map( A => mult_42_I5_n67, ZN => 
                           mult_42_I5_n304);
   mult_42_I5_U56 : HA_X1 port map( A => mult_42_I5_n148, B => mult_42_I5_n157,
                           CO => mult_42_I5_n89, S => mult_42_I5_n90);
   mult_42_I5_U55 : FA_X1 port map( A => mult_42_I5_n156, B => mult_42_I5_n139,
                           CI => mult_42_I5_n147, CO => mult_42_I5_n87, S => 
                           mult_42_I5_n88);
   mult_42_I5_U54 : HA_X1 port map( A => mult_42_I5_n107, B => mult_42_I5_n138,
                           CO => mult_42_I5_n85, S => mult_42_I5_n86);
   mult_42_I5_U53 : FA_X1 port map( A => mult_42_I5_n146, B => mult_42_I5_n155,
                           CI => mult_42_I5_n86, CO => mult_42_I5_n83, S => 
                           mult_42_I5_n84);
   mult_42_I5_U52 : FA_X1 port map( A => mult_42_I5_n154, B => mult_42_I5_n129,
                           CI => mult_42_I5_n145, CO => mult_42_I5_n81, S => 
                           mult_42_I5_n82);
   mult_42_I5_U51 : FA_X1 port map( A => mult_42_I5_n85, B => mult_42_I5_n137, 
                           CI => mult_42_I5_n82, CO => mult_42_I5_n79, S => 
                           mult_42_I5_n80);
   mult_42_I5_U50 : HA_X1 port map( A => mult_42_I5_n106, B => mult_42_I5_n128,
                           CO => mult_42_I5_n77, S => mult_42_I5_n78);
   mult_42_I5_U49 : FA_X1 port map( A => mult_42_I5_n136, B => mult_42_I5_n153,
                           CI => mult_42_I5_n144, CO => mult_42_I5_n75, S => 
                           mult_42_I5_n76);
   mult_42_I5_U48 : FA_X1 port map( A => mult_42_I5_n81, B => mult_42_I5_n78, 
                           CI => mult_42_I5_n76, CO => mult_42_I5_n73, S => 
                           mult_42_I5_n74);
   mult_42_I5_U47 : FA_X1 port map( A => mult_42_I5_n135, B => mult_42_I5_n119,
                           CI => mult_42_I5_n152, CO => mult_42_I5_n71, S => 
                           mult_42_I5_n72);
   mult_42_I5_U46 : FA_X1 port map( A => mult_42_I5_n127, B => mult_42_I5_n143,
                           CI => mult_42_I5_n77, CO => mult_42_I5_n69, S => 
                           mult_42_I5_n70);
   mult_42_I5_U45 : FA_X1 port map( A => mult_42_I5_n72, B => mult_42_I5_n75, 
                           CI => mult_42_I5_n70, CO => mult_42_I5_n67, S => 
                           mult_42_I5_n68);
   mult_42_I5_U44 : HA_X1 port map( A => mult_42_I5_n105, B => mult_42_I5_n118,
                           CO => mult_42_I5_n65, S => mult_42_I5_n66);
   mult_42_I5_U43 : FA_X1 port map( A => mult_42_I5_n126, B => mult_42_I5_n134,
                           CI => mult_42_I5_n142, CO => mult_42_I5_n63, S => 
                           mult_42_I5_n64);
   mult_42_I5_U42 : FA_X1 port map( A => mult_42_I5_n66, B => mult_42_I5_n151, 
                           CI => mult_42_I5_n71, CO => mult_42_I5_n61, S => 
                           mult_42_I5_n62);
   mult_42_I5_U41 : FA_X1 port map( A => mult_42_I5_n64, B => mult_42_I5_n69, 
                           CI => mult_42_I5_n62, CO => mult_42_I5_n59, S => 
                           mult_42_I5_n60);
   mult_42_I5_U38 : FA_X1 port map( A => mult_42_I5_n133, B => mult_42_I5_n117,
                           CI => mult_42_I5_n295, CO => mult_42_I5_n55, S => 
                           mult_42_I5_n56);
   mult_42_I5_U37 : FA_X1 port map( A => mult_42_I5_n58, B => mult_42_I5_n65, 
                           CI => mult_42_I5_n63, CO => mult_42_I5_n53, S => 
                           mult_42_I5_n54);
   mult_42_I5_U36 : FA_X1 port map( A => mult_42_I5_n61, B => mult_42_I5_n56, 
                           CI => mult_42_I5_n54, CO => mult_42_I5_n51, S => 
                           mult_42_I5_n52);
   mult_42_I5_U34 : FA_X1 port map( A => mult_42_I5_n124, B => mult_42_I5_n116,
                           CI => mult_42_I5_n132, CO => mult_42_I5_n47, S => 
                           mult_42_I5_n48);
   mult_42_I5_U33 : FA_X1 port map( A => mult_42_I5_n57, B => mult_42_I5_n50, 
                           CI => mult_42_I5_n55, CO => mult_42_I5_n45, S => 
                           mult_42_I5_n46);
   mult_42_I5_U32 : FA_X1 port map( A => mult_42_I5_n53, B => mult_42_I5_n48, 
                           CI => mult_42_I5_n46, CO => mult_42_I5_n43, S => 
                           mult_42_I5_n44);
   mult_42_I5_U31 : FA_X1 port map( A => mult_42_I5_n123, B => mult_42_I5_n115,
                           CI => mult_42_I5_n140, CO => mult_42_I5_n41, S => 
                           mult_42_I5_n42);
   mult_42_I5_U30 : FA_X1 port map( A => mult_42_I5_n297, B => mult_42_I5_n131,
                           CI => mult_42_I5_n47, CO => mult_42_I5_n39, S => 
                           mult_42_I5_n40);
   mult_42_I5_U29 : FA_X1 port map( A => mult_42_I5_n45, B => mult_42_I5_n42, 
                           CI => mult_42_I5_n40, CO => mult_42_I5_n37, S => 
                           mult_42_I5_n38);
   mult_42_I5_U27 : FA_X1 port map( A => mult_42_I5_n114, B => mult_42_I5_n122,
                           CI => mult_42_I5_n299, CO => mult_42_I5_n33, S => 
                           mult_42_I5_n34);
   mult_42_I5_U26 : FA_X1 port map( A => mult_42_I5_n34, B => mult_42_I5_n41, 
                           CI => mult_42_I5_n39, CO => mult_42_I5_n31, S => 
                           mult_42_I5_n32);
   mult_42_I5_U25 : FA_X1 port map( A => mult_42_I5_n121, B => mult_42_I5_n35, 
                           CI => mult_42_I5_n298, CO => mult_42_I5_n29, S => 
                           mult_42_I5_n30);
   mult_42_I5_U24 : FA_X1 port map( A => mult_42_I5_n33, B => mult_42_I5_n113, 
                           CI => mult_42_I5_n30, CO => mult_42_I5_n27, S => 
                           mult_42_I5_n28);
   mult_42_I5_U22 : FA_X1 port map( A => mult_42_I5_n301, B => mult_42_I5_n112,
                           CI => mult_42_I5_n29, CO => mult_42_I5_n23, S => 
                           mult_42_I5_n24);
   mult_42_I5_U21 : FA_X1 port map( A => mult_42_I5_n111, B => mult_42_I5_n25, 
                           CI => mult_42_I5_n300, CO => mult_42_I5_n21, S => 
                           mult_42_I5_n22);
   mult_42_I5_U10 : FA_X1 port map( A => mult_42_I5_n52, B => mult_42_I5_n59, 
                           CI => mult_42_I5_n10, CO => mult_42_I5_n9, S => N73)
                           ;
   mult_42_I5_U9 : FA_X1 port map( A => mult_42_I5_n44, B => mult_42_I5_n51, CI
                           => mult_42_I5_n9, CO => mult_42_I5_n8, S => N74);
   mult_42_I5_U8 : FA_X1 port map( A => mult_42_I5_n38, B => mult_42_I5_n43, CI
                           => mult_42_I5_n8, CO => mult_42_I5_n7, S => N75);
   mult_42_I5_U7 : FA_X1 port map( A => mult_42_I5_n32, B => mult_42_I5_n37, CI
                           => mult_42_I5_n7, CO => mult_42_I5_n6, S => N76);
   mult_42_I5_U6 : FA_X1 port map( A => mult_42_I5_n28, B => mult_42_I5_n31, CI
                           => mult_42_I5_n6, CO => mult_42_I5_n5, S => N77);
   mult_42_I5_U5 : FA_X1 port map( A => mult_42_I5_n24, B => mult_42_I5_n27, CI
                           => mult_42_I5_n5, CO => mult_42_I5_n4, S => N78);
   mult_42_I5_U4 : FA_X1 port map( A => mult_42_I5_n23, B => mult_42_I5_n22, CI
                           => mult_42_I5_n4, CO => mult_42_I5_n3, S => N79);
   mult_42_I5_U3 : FA_X1 port map( A => mult_42_I5_n21, B => mult_42_I5_n303, 
                           CI => mult_42_I5_n3, CO => mult_42_I5_n2, S => N80);
   mult_42_I5_U2 : FA_X1 port map( A => mult_42_I5_n302, B => mult_42_I5_n19, 
                           CI => mult_42_I5_n2, CO => mult_42_I5_n1, S => N81);
   mult_42_I6_U391 : NAND2_X1 port map( A1 => x_vector_51_port, A2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n341);
   mult_42_I6_U390 : XNOR2_X1 port map( A => B(52), B => x_vector_51_port, ZN 
                           => mult_42_I6_n340);
   mult_42_I6_U389 : OAI22_X1 port map( A1 => B(51), A2 => mult_42_I6_n341, B1 
                           => mult_42_I6_n340, B2 => mult_42_I6_n320, ZN => 
                           mult_42_I6_n402);
   mult_42_I6_U388 : NAND3_X1 port map( A1 => mult_42_I6_n402, A2 => 
                           mult_42_I6_n312, A3 => x_vector_51_port, ZN => 
                           mult_42_I6_n400);
   mult_42_I6_U387 : XNOR2_X1 port map( A => x_vector_52_port, B => 
                           x_vector_51_port, ZN => mult_42_I6_n352);
   mult_42_I6_U386 : NAND2_X1 port map( A1 => mult_42_I6_n319, A2 => 
                           mult_42_I6_n402, ZN => mult_42_I6_n401);
   mult_42_I6_U385 : MUX2_X1 port map( A => mult_42_I6_n400, B => 
                           mult_42_I6_n401, S => B(50), Z => mult_42_I6_n396);
   mult_42_I6_U384 : XOR2_X1 port map( A => x_vector_53_port, B => 
                           x_vector_52_port, Z => mult_42_I6_n399);
   mult_42_I6_U383 : NAND2_X1 port map( A1 => mult_42_I6_n352, A2 => 
                           mult_42_I6_n399, ZN => mult_42_I6_n351);
   mult_42_I6_U382 : NOR3_X1 port map( A1 => mult_42_I6_n352, A2 => B(50), A3 
                           => mult_42_I6_n317, ZN => mult_42_I6_n398);
   mult_42_I6_U381 : AOI21_X1 port map( B1 => x_vector_53_port, B2 => 
                           mult_42_I6_n318, A => mult_42_I6_n398, ZN => 
                           mult_42_I6_n397);
   mult_42_I6_U380 : OAI222_X1 port map( A1 => mult_42_I6_n396, A2 => 
                           mult_42_I6_n311, B1 => mult_42_I6_n397, B2 => 
                           mult_42_I6_n396, C1 => mult_42_I6_n397, C2 => 
                           mult_42_I6_n311, ZN => mult_42_I6_n395);
   mult_42_I6_U379 : AOI222_X1 port map( A1 => mult_42_I6_n395, A2 => 
                           mult_42_I6_n88, B1 => mult_42_I6_n395, B2 => 
                           mult_42_I6_n89, C1 => mult_42_I6_n89, C2 => 
                           mult_42_I6_n88, ZN => mult_42_I6_n394);
   mult_42_I6_U378 : OAI222_X1 port map( A1 => mult_42_I6_n394, A2 => 
                           mult_42_I6_n308, B1 => mult_42_I6_n394, B2 => 
                           mult_42_I6_n309, C1 => mult_42_I6_n309, C2 => 
                           mult_42_I6_n308, ZN => mult_42_I6_n393);
   mult_42_I6_U377 : AOI222_X1 port map( A1 => mult_42_I6_n393, A2 => 
                           mult_42_I6_n80, B1 => mult_42_I6_n393, B2 => 
                           mult_42_I6_n83, C1 => mult_42_I6_n83, C2 => 
                           mult_42_I6_n80, ZN => mult_42_I6_n392);
   mult_42_I6_U376 : OAI222_X1 port map( A1 => mult_42_I6_n392, A2 => 
                           mult_42_I6_n305, B1 => mult_42_I6_n392, B2 => 
                           mult_42_I6_n307, C1 => mult_42_I6_n307, C2 => 
                           mult_42_I6_n305, ZN => mult_42_I6_n391);
   mult_42_I6_U375 : AOI222_X1 port map( A1 => mult_42_I6_n391, A2 => 
                           mult_42_I6_n68, B1 => mult_42_I6_n391, B2 => 
                           mult_42_I6_n73, C1 => mult_42_I6_n73, C2 => 
                           mult_42_I6_n68, ZN => mult_42_I6_n390);
   mult_42_I6_U374 : OAI222_X1 port map( A1 => mult_42_I6_n390, A2 => 
                           mult_42_I6_n296, B1 => mult_42_I6_n390, B2 => 
                           mult_42_I6_n304, C1 => mult_42_I6_n304, C2 => 
                           mult_42_I6_n296, ZN => mult_42_I6_n10);
   mult_42_I6_U373 : XOR2_X1 port map( A => x_vector_59_port, B => 
                           x_vector_58_port, Z => mult_42_I6_n389);
   mult_42_I6_U372 : NAND2_X1 port map( A1 => mult_42_I6_n338, A2 => 
                           mult_42_I6_n389, ZN => mult_42_I6_n337);
   mult_42_I6_U371 : OR3_X1 port map( A1 => mult_42_I6_n338, A2 => B(50), A3 =>
                           mult_42_I6_n314, ZN => mult_42_I6_n388);
   mult_42_I6_U370 : OAI21_X1 port map( B1 => mult_42_I6_n314, B2 => 
                           mult_42_I6_n337, A => mult_42_I6_n388, ZN => 
                           mult_42_I6_n105);
   mult_42_I6_U369 : XOR2_X1 port map( A => x_vector_57_port, B => 
                           x_vector_56_port, Z => mult_42_I6_n387);
   mult_42_I6_U368 : NAND2_X1 port map( A1 => mult_42_I6_n327, A2 => 
                           mult_42_I6_n387, ZN => mult_42_I6_n326);
   mult_42_I6_U367 : OR3_X1 port map( A1 => mult_42_I6_n327, A2 => B(50), A3 =>
                           mult_42_I6_n315, ZN => mult_42_I6_n386);
   mult_42_I6_U366 : OAI21_X1 port map( B1 => mult_42_I6_n315, B2 => 
                           mult_42_I6_n326, A => mult_42_I6_n386, ZN => 
                           mult_42_I6_n106);
   mult_42_I6_U365 : XOR2_X1 port map( A => x_vector_55_port, B => 
                           x_vector_54_port, Z => mult_42_I6_n385);
   mult_42_I6_U364 : NAND2_X1 port map( A1 => mult_42_I6_n332, A2 => 
                           mult_42_I6_n385, ZN => mult_42_I6_n331);
   mult_42_I6_U363 : OR3_X1 port map( A1 => mult_42_I6_n332, A2 => B(50), A3 =>
                           mult_42_I6_n316, ZN => mult_42_I6_n384);
   mult_42_I6_U362 : OAI21_X1 port map( B1 => mult_42_I6_n316, B2 => 
                           mult_42_I6_n331, A => mult_42_I6_n384, ZN => 
                           mult_42_I6_n107);
   mult_42_I6_U361 : XOR2_X1 port map( A => B(59), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n339);
   mult_42_I6_U360 : OAI22_X1 port map( A1 => mult_42_I6_n339, A2 => 
                           mult_42_I6_n338, B1 => mult_42_I6_n337, B2 => 
                           mult_42_I6_n339, ZN => mult_42_I6_n383);
   mult_42_I6_U359 : XOR2_X1 port map( A => B(57), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n382);
   mult_42_I6_U358 : XOR2_X1 port map( A => B(58), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n336);
   mult_42_I6_U357 : OAI22_X1 port map( A1 => mult_42_I6_n382, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n336, ZN => mult_42_I6_n111);
   mult_42_I6_U356 : XOR2_X1 port map( A => B(56), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n381);
   mult_42_I6_U355 : OAI22_X1 port map( A1 => mult_42_I6_n381, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n382, ZN => mult_42_I6_n112);
   mult_42_I6_U354 : XOR2_X1 port map( A => B(55), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n380);
   mult_42_I6_U353 : OAI22_X1 port map( A1 => mult_42_I6_n380, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n381, ZN => mult_42_I6_n113);
   mult_42_I6_U352 : XOR2_X1 port map( A => B(54), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n379);
   mult_42_I6_U351 : OAI22_X1 port map( A1 => mult_42_I6_n379, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n380, ZN => mult_42_I6_n114);
   mult_42_I6_U350 : XOR2_X1 port map( A => B(53), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n378);
   mult_42_I6_U349 : OAI22_X1 port map( A1 => mult_42_I6_n378, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n379, ZN => mult_42_I6_n115);
   mult_42_I6_U348 : XOR2_X1 port map( A => B(52), B => mult_42_I6_n314, Z => 
                           mult_42_I6_n377);
   mult_42_I6_U347 : OAI22_X1 port map( A1 => mult_42_I6_n377, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n378, ZN => mult_42_I6_n116);
   mult_42_I6_U346 : XOR2_X1 port map( A => mult_42_I6_n312, B => 
                           x_vector_59_port, Z => mult_42_I6_n376);
   mult_42_I6_U345 : OAI22_X1 port map( A1 => mult_42_I6_n376, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n377, ZN => mult_42_I6_n117);
   mult_42_I6_U344 : XOR2_X1 port map( A => mult_42_I6_n314, B => B(50), Z => 
                           mult_42_I6_n375);
   mult_42_I6_U343 : OAI22_X1 port map( A1 => mult_42_I6_n375, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n376, ZN => mult_42_I6_n118);
   mult_42_I6_U342 : NOR2_X1 port map( A1 => mult_42_I6_n338, A2 => 
                           mult_42_I6_n313, ZN => mult_42_I6_n119);
   mult_42_I6_U341 : XOR2_X1 port map( A => B(59), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n335);
   mult_42_I6_U340 : OAI22_X1 port map( A1 => mult_42_I6_n335, A2 => 
                           mult_42_I6_n327, B1 => mult_42_I6_n326, B2 => 
                           mult_42_I6_n335, ZN => mult_42_I6_n374);
   mult_42_I6_U339 : XOR2_X1 port map( A => B(57), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n373);
   mult_42_I6_U338 : XOR2_X1 port map( A => B(58), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n334);
   mult_42_I6_U337 : OAI22_X1 port map( A1 => mult_42_I6_n373, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n334, ZN => mult_42_I6_n121);
   mult_42_I6_U336 : XOR2_X1 port map( A => B(56), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n372);
   mult_42_I6_U335 : OAI22_X1 port map( A1 => mult_42_I6_n372, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n373, ZN => mult_42_I6_n122);
   mult_42_I6_U334 : XOR2_X1 port map( A => B(55), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n371);
   mult_42_I6_U333 : OAI22_X1 port map( A1 => mult_42_I6_n371, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n372, ZN => mult_42_I6_n123);
   mult_42_I6_U332 : XOR2_X1 port map( A => B(54), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n328);
   mult_42_I6_U331 : OAI22_X1 port map( A1 => mult_42_I6_n328, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n371, ZN => mult_42_I6_n124);
   mult_42_I6_U330 : XOR2_X1 port map( A => B(52), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n370);
   mult_42_I6_U329 : XOR2_X1 port map( A => B(53), B => mult_42_I6_n315, Z => 
                           mult_42_I6_n325);
   mult_42_I6_U328 : OAI22_X1 port map( A1 => mult_42_I6_n370, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n325, ZN => mult_42_I6_n126);
   mult_42_I6_U327 : XOR2_X1 port map( A => mult_42_I6_n312, B => 
                           x_vector_57_port, Z => mult_42_I6_n369);
   mult_42_I6_U326 : OAI22_X1 port map( A1 => mult_42_I6_n369, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n370, ZN => mult_42_I6_n127);
   mult_42_I6_U325 : XOR2_X1 port map( A => mult_42_I6_n313, B => 
                           x_vector_57_port, Z => mult_42_I6_n368);
   mult_42_I6_U324 : OAI22_X1 port map( A1 => mult_42_I6_n368, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n369, ZN => mult_42_I6_n128);
   mult_42_I6_U323 : NOR2_X1 port map( A1 => mult_42_I6_n327, A2 => 
                           mult_42_I6_n313, ZN => mult_42_I6_n129);
   mult_42_I6_U322 : XOR2_X1 port map( A => B(59), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n333);
   mult_42_I6_U321 : OAI22_X1 port map( A1 => mult_42_I6_n333, A2 => 
                           mult_42_I6_n332, B1 => mult_42_I6_n331, B2 => 
                           mult_42_I6_n333, ZN => mult_42_I6_n367);
   mult_42_I6_U320 : XOR2_X1 port map( A => B(57), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n366);
   mult_42_I6_U319 : XOR2_X1 port map( A => B(58), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n330);
   mult_42_I6_U318 : OAI22_X1 port map( A1 => mult_42_I6_n366, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n330, ZN => mult_42_I6_n131);
   mult_42_I6_U317 : XOR2_X1 port map( A => B(56), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n365);
   mult_42_I6_U316 : OAI22_X1 port map( A1 => mult_42_I6_n365, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n366, ZN => mult_42_I6_n132);
   mult_42_I6_U315 : XOR2_X1 port map( A => B(55), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n364);
   mult_42_I6_U314 : OAI22_X1 port map( A1 => mult_42_I6_n364, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n365, ZN => mult_42_I6_n133);
   mult_42_I6_U313 : XOR2_X1 port map( A => B(54), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n363);
   mult_42_I6_U312 : OAI22_X1 port map( A1 => mult_42_I6_n363, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n364, ZN => mult_42_I6_n134);
   mult_42_I6_U311 : XOR2_X1 port map( A => B(53), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n362);
   mult_42_I6_U310 : OAI22_X1 port map( A1 => mult_42_I6_n362, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n363, ZN => mult_42_I6_n135);
   mult_42_I6_U309 : XOR2_X1 port map( A => B(52), B => mult_42_I6_n316, Z => 
                           mult_42_I6_n361);
   mult_42_I6_U308 : OAI22_X1 port map( A1 => mult_42_I6_n361, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n362, ZN => mult_42_I6_n136);
   mult_42_I6_U307 : XOR2_X1 port map( A => mult_42_I6_n312, B => 
                           x_vector_55_port, Z => mult_42_I6_n360);
   mult_42_I6_U306 : OAI22_X1 port map( A1 => mult_42_I6_n360, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n361, ZN => mult_42_I6_n137);
   mult_42_I6_U305 : XOR2_X1 port map( A => mult_42_I6_n313, B => 
                           x_vector_55_port, Z => mult_42_I6_n359);
   mult_42_I6_U304 : OAI22_X1 port map( A1 => mult_42_I6_n359, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n360, ZN => mult_42_I6_n138);
   mult_42_I6_U303 : NOR2_X1 port map( A1 => mult_42_I6_n332, A2 => 
                           mult_42_I6_n313, ZN => mult_42_I6_n139);
   mult_42_I6_U302 : XOR2_X1 port map( A => B(59), B => x_vector_53_port, Z => 
                           mult_42_I6_n329);
   mult_42_I6_U301 : AOI22_X1 port map( A1 => mult_42_I6_n329, A2 => 
                           mult_42_I6_n319, B1 => mult_42_I6_n318, B2 => 
                           mult_42_I6_n329, ZN => mult_42_I6_n140);
   mult_42_I6_U300 : XOR2_X1 port map( A => B(56), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n358);
   mult_42_I6_U299 : XOR2_X1 port map( A => B(57), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n324);
   mult_42_I6_U298 : OAI22_X1 port map( A1 => mult_42_I6_n358, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n324, ZN => mult_42_I6_n142);
   mult_42_I6_U297 : XOR2_X1 port map( A => B(55), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n357);
   mult_42_I6_U296 : OAI22_X1 port map( A1 => mult_42_I6_n357, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n358, ZN => mult_42_I6_n143);
   mult_42_I6_U295 : XOR2_X1 port map( A => B(54), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n356);
   mult_42_I6_U294 : OAI22_X1 port map( A1 => mult_42_I6_n356, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n357, ZN => mult_42_I6_n144);
   mult_42_I6_U293 : XOR2_X1 port map( A => B(53), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n355);
   mult_42_I6_U292 : OAI22_X1 port map( A1 => mult_42_I6_n355, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n356, ZN => mult_42_I6_n145);
   mult_42_I6_U291 : XOR2_X1 port map( A => B(52), B => mult_42_I6_n317, Z => 
                           mult_42_I6_n354);
   mult_42_I6_U290 : OAI22_X1 port map( A1 => mult_42_I6_n354, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n355, ZN => mult_42_I6_n146);
   mult_42_I6_U289 : XOR2_X1 port map( A => mult_42_I6_n312, B => 
                           x_vector_53_port, Z => mult_42_I6_n353);
   mult_42_I6_U288 : OAI22_X1 port map( A1 => mult_42_I6_n353, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n354, ZN => mult_42_I6_n147);
   mult_42_I6_U287 : XOR2_X1 port map( A => mult_42_I6_n313, B => 
                           x_vector_53_port, Z => mult_42_I6_n350);
   mult_42_I6_U286 : OAI22_X1 port map( A1 => mult_42_I6_n350, A2 => 
                           mult_42_I6_n351, B1 => mult_42_I6_n352, B2 => 
                           mult_42_I6_n353, ZN => mult_42_I6_n148);
   mult_42_I6_U285 : XNOR2_X1 port map( A => B(59), B => x_vector_51_port, ZN 
                           => mult_42_I6_n348);
   mult_42_I6_U284 : OAI22_X1 port map( A1 => mult_42_I6_n320, A2 => 
                           mult_42_I6_n348, B1 => mult_42_I6_n341, B2 => 
                           mult_42_I6_n348, ZN => mult_42_I6_n349);
   mult_42_I6_U283 : XNOR2_X1 port map( A => B(58), B => x_vector_51_port, ZN 
                           => mult_42_I6_n347);
   mult_42_I6_U282 : OAI22_X1 port map( A1 => mult_42_I6_n347, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n348, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n151);
   mult_42_I6_U281 : XNOR2_X1 port map( A => B(57), B => x_vector_51_port, ZN 
                           => mult_42_I6_n346);
   mult_42_I6_U280 : OAI22_X1 port map( A1 => mult_42_I6_n346, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n347, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n152);
   mult_42_I6_U279 : XNOR2_X1 port map( A => B(56), B => x_vector_51_port, ZN 
                           => mult_42_I6_n345);
   mult_42_I6_U278 : OAI22_X1 port map( A1 => mult_42_I6_n345, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n346, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n153);
   mult_42_I6_U277 : XNOR2_X1 port map( A => B(55), B => x_vector_51_port, ZN 
                           => mult_42_I6_n344);
   mult_42_I6_U276 : OAI22_X1 port map( A1 => mult_42_I6_n344, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n345, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n154);
   mult_42_I6_U275 : XNOR2_X1 port map( A => B(54), B => x_vector_51_port, ZN 
                           => mult_42_I6_n343);
   mult_42_I6_U274 : OAI22_X1 port map( A1 => mult_42_I6_n343, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n344, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n155);
   mult_42_I6_U273 : XNOR2_X1 port map( A => B(53), B => x_vector_51_port, ZN 
                           => mult_42_I6_n342);
   mult_42_I6_U272 : OAI22_X1 port map( A1 => mult_42_I6_n342, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n343, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n156);
   mult_42_I6_U271 : OAI22_X1 port map( A1 => mult_42_I6_n340, A2 => 
                           mult_42_I6_n341, B1 => mult_42_I6_n342, B2 => 
                           mult_42_I6_n320, ZN => mult_42_I6_n157);
   mult_42_I6_U270 : OAI22_X1 port map( A1 => mult_42_I6_n336, A2 => 
                           mult_42_I6_n337, B1 => mult_42_I6_n338, B2 => 
                           mult_42_I6_n339, ZN => mult_42_I6_n19);
   mult_42_I6_U269 : OAI22_X1 port map( A1 => mult_42_I6_n334, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n335, ZN => mult_42_I6_n25);
   mult_42_I6_U268 : OAI22_X1 port map( A1 => mult_42_I6_n330, A2 => 
                           mult_42_I6_n331, B1 => mult_42_I6_n332, B2 => 
                           mult_42_I6_n333, ZN => mult_42_I6_n35);
   mult_42_I6_U267 : XOR2_X1 port map( A => B(58), B => x_vector_53_port, Z => 
                           mult_42_I6_n323);
   mult_42_I6_U266 : AOI22_X1 port map( A1 => mult_42_I6_n323, A2 => 
                           mult_42_I6_n318, B1 => mult_42_I6_n319, B2 => 
                           mult_42_I6_n329, ZN => mult_42_I6_n50);
   mult_42_I6_U265 : OAI22_X1 port map( A1 => mult_42_I6_n325, A2 => 
                           mult_42_I6_n326, B1 => mult_42_I6_n327, B2 => 
                           mult_42_I6_n328, ZN => mult_42_I6_n321);
   mult_42_I6_U264 : AOI22_X1 port map( A1 => mult_42_I6_n306, A2 => 
                           mult_42_I6_n318, B1 => mult_42_I6_n319, B2 => 
                           mult_42_I6_n323, ZN => mult_42_I6_n322);
   mult_42_I6_U263 : NAND2_X1 port map( A1 => mult_42_I6_n310, A2 => 
                           mult_42_I6_n322, ZN => mult_42_I6_n57);
   mult_42_I6_U262 : XOR2_X1 port map( A => mult_42_I6_n321, B => 
                           mult_42_I6_n322, Z => mult_42_I6_n58);
   mult_42_I6_U261 : XNOR2_X2 port map( A => x_vector_58_port, B => 
                           x_vector_57_port, ZN => mult_42_I6_n338);
   mult_42_I6_U260 : XNOR2_X2 port map( A => x_vector_56_port, B => 
                           x_vector_55_port, ZN => mult_42_I6_n327);
   mult_42_I6_U259 : XNOR2_X2 port map( A => x_vector_54_port, B => 
                           x_vector_53_port, ZN => mult_42_I6_n332);
   mult_42_I6_U258 : INV_X1 port map( A => B(51), ZN => mult_42_I6_n312);
   mult_42_I6_U257 : INV_X1 port map( A => B(50), ZN => mult_42_I6_n313);
   mult_42_I6_U256 : INV_X1 port map( A => x_vector_53_port, ZN => 
                           mult_42_I6_n317);
   mult_42_I6_U255 : INV_X1 port map( A => x_vector_50_port, ZN => 
                           mult_42_I6_n320);
   mult_42_I6_U254 : INV_X1 port map( A => x_vector_57_port, ZN => 
                           mult_42_I6_n315);
   mult_42_I6_U253 : INV_X1 port map( A => x_vector_55_port, ZN => 
                           mult_42_I6_n316);
   mult_42_I6_U252 : INV_X1 port map( A => x_vector_59_port, ZN => 
                           mult_42_I6_n314);
   mult_42_I6_U251 : INV_X1 port map( A => mult_42_I6_n367, ZN => 
                           mult_42_I6_n298);
   mult_42_I6_U250 : INV_X1 port map( A => mult_42_I6_n374, ZN => 
                           mult_42_I6_n300);
   mult_42_I6_U249 : INV_X1 port map( A => mult_42_I6_n25, ZN => 
                           mult_42_I6_n301);
   mult_42_I6_U248 : INV_X1 port map( A => mult_42_I6_n35, ZN => 
                           mult_42_I6_n299);
   mult_42_I6_U247 : INV_X1 port map( A => mult_42_I6_n90, ZN => 
                           mult_42_I6_n311);
   mult_42_I6_U246 : INV_X1 port map( A => mult_42_I6_n50, ZN => 
                           mult_42_I6_n297);
   mult_42_I6_U245 : INV_X1 port map( A => mult_42_I6_n349, ZN => 
                           mult_42_I6_n295);
   mult_42_I6_U244 : INV_X1 port map( A => mult_42_I6_n383, ZN => 
                           mult_42_I6_n302);
   mult_42_I6_U243 : INV_X1 port map( A => mult_42_I6_n351, ZN => 
                           mult_42_I6_n318);
   mult_42_I6_U242 : INV_X1 port map( A => mult_42_I6_n352, ZN => 
                           mult_42_I6_n319);
   mult_42_I6_U241 : INV_X1 port map( A => mult_42_I6_n324, ZN => 
                           mult_42_I6_n306);
   mult_42_I6_U240 : INV_X1 port map( A => mult_42_I6_n84, ZN => 
                           mult_42_I6_n308);
   mult_42_I6_U239 : INV_X1 port map( A => mult_42_I6_n87, ZN => 
                           mult_42_I6_n309);
   mult_42_I6_U238 : INV_X1 port map( A => mult_42_I6_n19, ZN => 
                           mult_42_I6_n303);
   mult_42_I6_U237 : INV_X1 port map( A => mult_42_I6_n321, ZN => 
                           mult_42_I6_n310);
   mult_42_I6_U236 : INV_X1 port map( A => mult_42_I6_n1, ZN => N102);
   mult_42_I6_U235 : INV_X1 port map( A => mult_42_I6_n74, ZN => 
                           mult_42_I6_n305);
   mult_42_I6_U234 : INV_X1 port map( A => mult_42_I6_n79, ZN => 
                           mult_42_I6_n307);
   mult_42_I6_U233 : INV_X1 port map( A => mult_42_I6_n60, ZN => 
                           mult_42_I6_n296);
   mult_42_I6_U232 : INV_X1 port map( A => mult_42_I6_n67, ZN => 
                           mult_42_I6_n304);
   mult_42_I6_U56 : HA_X1 port map( A => mult_42_I6_n148, B => mult_42_I6_n157,
                           CO => mult_42_I6_n89, S => mult_42_I6_n90);
   mult_42_I6_U55 : FA_X1 port map( A => mult_42_I6_n156, B => mult_42_I6_n139,
                           CI => mult_42_I6_n147, CO => mult_42_I6_n87, S => 
                           mult_42_I6_n88);
   mult_42_I6_U54 : HA_X1 port map( A => mult_42_I6_n107, B => mult_42_I6_n138,
                           CO => mult_42_I6_n85, S => mult_42_I6_n86);
   mult_42_I6_U53 : FA_X1 port map( A => mult_42_I6_n146, B => mult_42_I6_n155,
                           CI => mult_42_I6_n86, CO => mult_42_I6_n83, S => 
                           mult_42_I6_n84);
   mult_42_I6_U52 : FA_X1 port map( A => mult_42_I6_n154, B => mult_42_I6_n129,
                           CI => mult_42_I6_n145, CO => mult_42_I6_n81, S => 
                           mult_42_I6_n82);
   mult_42_I6_U51 : FA_X1 port map( A => mult_42_I6_n85, B => mult_42_I6_n137, 
                           CI => mult_42_I6_n82, CO => mult_42_I6_n79, S => 
                           mult_42_I6_n80);
   mult_42_I6_U50 : HA_X1 port map( A => mult_42_I6_n106, B => mult_42_I6_n128,
                           CO => mult_42_I6_n77, S => mult_42_I6_n78);
   mult_42_I6_U49 : FA_X1 port map( A => mult_42_I6_n136, B => mult_42_I6_n153,
                           CI => mult_42_I6_n144, CO => mult_42_I6_n75, S => 
                           mult_42_I6_n76);
   mult_42_I6_U48 : FA_X1 port map( A => mult_42_I6_n81, B => mult_42_I6_n78, 
                           CI => mult_42_I6_n76, CO => mult_42_I6_n73, S => 
                           mult_42_I6_n74);
   mult_42_I6_U47 : FA_X1 port map( A => mult_42_I6_n135, B => mult_42_I6_n119,
                           CI => mult_42_I6_n152, CO => mult_42_I6_n71, S => 
                           mult_42_I6_n72);
   mult_42_I6_U46 : FA_X1 port map( A => mult_42_I6_n127, B => mult_42_I6_n143,
                           CI => mult_42_I6_n77, CO => mult_42_I6_n69, S => 
                           mult_42_I6_n70);
   mult_42_I6_U45 : FA_X1 port map( A => mult_42_I6_n72, B => mult_42_I6_n75, 
                           CI => mult_42_I6_n70, CO => mult_42_I6_n67, S => 
                           mult_42_I6_n68);
   mult_42_I6_U44 : HA_X1 port map( A => mult_42_I6_n105, B => mult_42_I6_n118,
                           CO => mult_42_I6_n65, S => mult_42_I6_n66);
   mult_42_I6_U43 : FA_X1 port map( A => mult_42_I6_n126, B => mult_42_I6_n134,
                           CI => mult_42_I6_n142, CO => mult_42_I6_n63, S => 
                           mult_42_I6_n64);
   mult_42_I6_U42 : FA_X1 port map( A => mult_42_I6_n66, B => mult_42_I6_n151, 
                           CI => mult_42_I6_n71, CO => mult_42_I6_n61, S => 
                           mult_42_I6_n62);
   mult_42_I6_U41 : FA_X1 port map( A => mult_42_I6_n64, B => mult_42_I6_n69, 
                           CI => mult_42_I6_n62, CO => mult_42_I6_n59, S => 
                           mult_42_I6_n60);
   mult_42_I6_U38 : FA_X1 port map( A => mult_42_I6_n133, B => mult_42_I6_n117,
                           CI => mult_42_I6_n295, CO => mult_42_I6_n55, S => 
                           mult_42_I6_n56);
   mult_42_I6_U37 : FA_X1 port map( A => mult_42_I6_n58, B => mult_42_I6_n65, 
                           CI => mult_42_I6_n63, CO => mult_42_I6_n53, S => 
                           mult_42_I6_n54);
   mult_42_I6_U36 : FA_X1 port map( A => mult_42_I6_n61, B => mult_42_I6_n56, 
                           CI => mult_42_I6_n54, CO => mult_42_I6_n51, S => 
                           mult_42_I6_n52);
   mult_42_I6_U34 : FA_X1 port map( A => mult_42_I6_n124, B => mult_42_I6_n116,
                           CI => mult_42_I6_n132, CO => mult_42_I6_n47, S => 
                           mult_42_I6_n48);
   mult_42_I6_U33 : FA_X1 port map( A => mult_42_I6_n57, B => mult_42_I6_n50, 
                           CI => mult_42_I6_n55, CO => mult_42_I6_n45, S => 
                           mult_42_I6_n46);
   mult_42_I6_U32 : FA_X1 port map( A => mult_42_I6_n53, B => mult_42_I6_n48, 
                           CI => mult_42_I6_n46, CO => mult_42_I6_n43, S => 
                           mult_42_I6_n44);
   mult_42_I6_U31 : FA_X1 port map( A => mult_42_I6_n123, B => mult_42_I6_n115,
                           CI => mult_42_I6_n140, CO => mult_42_I6_n41, S => 
                           mult_42_I6_n42);
   mult_42_I6_U30 : FA_X1 port map( A => mult_42_I6_n297, B => mult_42_I6_n131,
                           CI => mult_42_I6_n47, CO => mult_42_I6_n39, S => 
                           mult_42_I6_n40);
   mult_42_I6_U29 : FA_X1 port map( A => mult_42_I6_n45, B => mult_42_I6_n42, 
                           CI => mult_42_I6_n40, CO => mult_42_I6_n37, S => 
                           mult_42_I6_n38);
   mult_42_I6_U27 : FA_X1 port map( A => mult_42_I6_n114, B => mult_42_I6_n122,
                           CI => mult_42_I6_n299, CO => mult_42_I6_n33, S => 
                           mult_42_I6_n34);
   mult_42_I6_U26 : FA_X1 port map( A => mult_42_I6_n34, B => mult_42_I6_n41, 
                           CI => mult_42_I6_n39, CO => mult_42_I6_n31, S => 
                           mult_42_I6_n32);
   mult_42_I6_U25 : FA_X1 port map( A => mult_42_I6_n121, B => mult_42_I6_n35, 
                           CI => mult_42_I6_n298, CO => mult_42_I6_n29, S => 
                           mult_42_I6_n30);
   mult_42_I6_U24 : FA_X1 port map( A => mult_42_I6_n33, B => mult_42_I6_n113, 
                           CI => mult_42_I6_n30, CO => mult_42_I6_n27, S => 
                           mult_42_I6_n28);
   mult_42_I6_U22 : FA_X1 port map( A => mult_42_I6_n301, B => mult_42_I6_n112,
                           CI => mult_42_I6_n29, CO => mult_42_I6_n23, S => 
                           mult_42_I6_n24);
   mult_42_I6_U21 : FA_X1 port map( A => mult_42_I6_n111, B => mult_42_I6_n25, 
                           CI => mult_42_I6_n300, CO => mult_42_I6_n21, S => 
                           mult_42_I6_n22);
   mult_42_I6_U10 : FA_X1 port map( A => mult_42_I6_n52, B => mult_42_I6_n59, 
                           CI => mult_42_I6_n10, CO => mult_42_I6_n9, S => N93)
                           ;
   mult_42_I6_U9 : FA_X1 port map( A => mult_42_I6_n44, B => mult_42_I6_n51, CI
                           => mult_42_I6_n9, CO => mult_42_I6_n8, S => N94);
   mult_42_I6_U8 : FA_X1 port map( A => mult_42_I6_n38, B => mult_42_I6_n43, CI
                           => mult_42_I6_n8, CO => mult_42_I6_n7, S => N95);
   mult_42_I6_U7 : FA_X1 port map( A => mult_42_I6_n32, B => mult_42_I6_n37, CI
                           => mult_42_I6_n7, CO => mult_42_I6_n6, S => N96);
   mult_42_I6_U6 : FA_X1 port map( A => mult_42_I6_n28, B => mult_42_I6_n31, CI
                           => mult_42_I6_n6, CO => mult_42_I6_n5, S => N97);
   mult_42_I6_U5 : FA_X1 port map( A => mult_42_I6_n24, B => mult_42_I6_n27, CI
                           => mult_42_I6_n5, CO => mult_42_I6_n4, S => N98);
   mult_42_I6_U4 : FA_X1 port map( A => mult_42_I6_n23, B => mult_42_I6_n22, CI
                           => mult_42_I6_n4, CO => mult_42_I6_n3, S => N99);
   mult_42_I6_U3 : FA_X1 port map( A => mult_42_I6_n21, B => mult_42_I6_n303, 
                           CI => mult_42_I6_n3, CO => mult_42_I6_n2, S => N100)
                           ;
   mult_42_I6_U2 : FA_X1 port map( A => mult_42_I6_n302, B => mult_42_I6_n19, 
                           CI => mult_42_I6_n2, CO => mult_42_I6_n1, S => N101)
                           ;
   mult_42_I7_U391 : NAND2_X1 port map( A1 => x_vector_61_port, A2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n341);
   mult_42_I7_U390 : XNOR2_X1 port map( A => B(62), B => x_vector_61_port, ZN 
                           => mult_42_I7_n340);
   mult_42_I7_U389 : OAI22_X1 port map( A1 => B(61), A2 => mult_42_I7_n341, B1 
                           => mult_42_I7_n340, B2 => mult_42_I7_n320, ZN => 
                           mult_42_I7_n402);
   mult_42_I7_U388 : NAND3_X1 port map( A1 => mult_42_I7_n402, A2 => 
                           mult_42_I7_n312, A3 => x_vector_61_port, ZN => 
                           mult_42_I7_n400);
   mult_42_I7_U387 : XNOR2_X1 port map( A => x_vector_62_port, B => 
                           x_vector_61_port, ZN => mult_42_I7_n352);
   mult_42_I7_U386 : NAND2_X1 port map( A1 => mult_42_I7_n319, A2 => 
                           mult_42_I7_n402, ZN => mult_42_I7_n401);
   mult_42_I7_U385 : MUX2_X1 port map( A => mult_42_I7_n400, B => 
                           mult_42_I7_n401, S => B(60), Z => mult_42_I7_n396);
   mult_42_I7_U384 : XOR2_X1 port map( A => x_vector_63_port, B => 
                           x_vector_62_port, Z => mult_42_I7_n399);
   mult_42_I7_U383 : NAND2_X1 port map( A1 => mult_42_I7_n352, A2 => 
                           mult_42_I7_n399, ZN => mult_42_I7_n351);
   mult_42_I7_U382 : NOR3_X1 port map( A1 => mult_42_I7_n352, A2 => B(60), A3 
                           => mult_42_I7_n317, ZN => mult_42_I7_n398);
   mult_42_I7_U381 : AOI21_X1 port map( B1 => x_vector_63_port, B2 => 
                           mult_42_I7_n318, A => mult_42_I7_n398, ZN => 
                           mult_42_I7_n397);
   mult_42_I7_U380 : OAI222_X1 port map( A1 => mult_42_I7_n396, A2 => 
                           mult_42_I7_n311, B1 => mult_42_I7_n397, B2 => 
                           mult_42_I7_n396, C1 => mult_42_I7_n397, C2 => 
                           mult_42_I7_n311, ZN => mult_42_I7_n395);
   mult_42_I7_U379 : AOI222_X1 port map( A1 => mult_42_I7_n395, A2 => 
                           mult_42_I7_n88, B1 => mult_42_I7_n395, B2 => 
                           mult_42_I7_n89, C1 => mult_42_I7_n89, C2 => 
                           mult_42_I7_n88, ZN => mult_42_I7_n394);
   mult_42_I7_U378 : OAI222_X1 port map( A1 => mult_42_I7_n394, A2 => 
                           mult_42_I7_n308, B1 => mult_42_I7_n394, B2 => 
                           mult_42_I7_n309, C1 => mult_42_I7_n309, C2 => 
                           mult_42_I7_n308, ZN => mult_42_I7_n393);
   mult_42_I7_U377 : AOI222_X1 port map( A1 => mult_42_I7_n393, A2 => 
                           mult_42_I7_n80, B1 => mult_42_I7_n393, B2 => 
                           mult_42_I7_n83, C1 => mult_42_I7_n83, C2 => 
                           mult_42_I7_n80, ZN => mult_42_I7_n392);
   mult_42_I7_U376 : OAI222_X1 port map( A1 => mult_42_I7_n392, A2 => 
                           mult_42_I7_n305, B1 => mult_42_I7_n392, B2 => 
                           mult_42_I7_n307, C1 => mult_42_I7_n307, C2 => 
                           mult_42_I7_n305, ZN => mult_42_I7_n391);
   mult_42_I7_U375 : AOI222_X1 port map( A1 => mult_42_I7_n391, A2 => 
                           mult_42_I7_n68, B1 => mult_42_I7_n391, B2 => 
                           mult_42_I7_n73, C1 => mult_42_I7_n73, C2 => 
                           mult_42_I7_n68, ZN => mult_42_I7_n390);
   mult_42_I7_U374 : OAI222_X1 port map( A1 => mult_42_I7_n390, A2 => 
                           mult_42_I7_n296, B1 => mult_42_I7_n390, B2 => 
                           mult_42_I7_n304, C1 => mult_42_I7_n304, C2 => 
                           mult_42_I7_n296, ZN => mult_42_I7_n10);
   mult_42_I7_U373 : XOR2_X1 port map( A => x_vector_69_port, B => 
                           x_vector_68_port, Z => mult_42_I7_n389);
   mult_42_I7_U372 : NAND2_X1 port map( A1 => mult_42_I7_n338, A2 => 
                           mult_42_I7_n389, ZN => mult_42_I7_n337);
   mult_42_I7_U371 : OR3_X1 port map( A1 => mult_42_I7_n338, A2 => B(60), A3 =>
                           mult_42_I7_n314, ZN => mult_42_I7_n388);
   mult_42_I7_U370 : OAI21_X1 port map( B1 => mult_42_I7_n314, B2 => 
                           mult_42_I7_n337, A => mult_42_I7_n388, ZN => 
                           mult_42_I7_n105);
   mult_42_I7_U369 : XOR2_X1 port map( A => x_vector_67_port, B => 
                           x_vector_66_port, Z => mult_42_I7_n387);
   mult_42_I7_U368 : NAND2_X1 port map( A1 => mult_42_I7_n327, A2 => 
                           mult_42_I7_n387, ZN => mult_42_I7_n326);
   mult_42_I7_U367 : OR3_X1 port map( A1 => mult_42_I7_n327, A2 => B(60), A3 =>
                           mult_42_I7_n315, ZN => mult_42_I7_n386);
   mult_42_I7_U366 : OAI21_X1 port map( B1 => mult_42_I7_n315, B2 => 
                           mult_42_I7_n326, A => mult_42_I7_n386, ZN => 
                           mult_42_I7_n106);
   mult_42_I7_U365 : XOR2_X1 port map( A => x_vector_65_port, B => 
                           x_vector_64_port, Z => mult_42_I7_n385);
   mult_42_I7_U364 : NAND2_X1 port map( A1 => mult_42_I7_n332, A2 => 
                           mult_42_I7_n385, ZN => mult_42_I7_n331);
   mult_42_I7_U363 : OR3_X1 port map( A1 => mult_42_I7_n332, A2 => B(60), A3 =>
                           mult_42_I7_n316, ZN => mult_42_I7_n384);
   mult_42_I7_U362 : OAI21_X1 port map( B1 => mult_42_I7_n316, B2 => 
                           mult_42_I7_n331, A => mult_42_I7_n384, ZN => 
                           mult_42_I7_n107);
   mult_42_I7_U361 : XOR2_X1 port map( A => B(69), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n339);
   mult_42_I7_U360 : OAI22_X1 port map( A1 => mult_42_I7_n339, A2 => 
                           mult_42_I7_n338, B1 => mult_42_I7_n337, B2 => 
                           mult_42_I7_n339, ZN => mult_42_I7_n383);
   mult_42_I7_U359 : XOR2_X1 port map( A => B(67), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n382);
   mult_42_I7_U358 : XOR2_X1 port map( A => B(68), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n336);
   mult_42_I7_U357 : OAI22_X1 port map( A1 => mult_42_I7_n382, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n336, ZN => mult_42_I7_n111);
   mult_42_I7_U356 : XOR2_X1 port map( A => B(66), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n381);
   mult_42_I7_U355 : OAI22_X1 port map( A1 => mult_42_I7_n381, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n382, ZN => mult_42_I7_n112);
   mult_42_I7_U354 : XOR2_X1 port map( A => B(65), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n380);
   mult_42_I7_U353 : OAI22_X1 port map( A1 => mult_42_I7_n380, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n381, ZN => mult_42_I7_n113);
   mult_42_I7_U352 : XOR2_X1 port map( A => B(64), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n379);
   mult_42_I7_U351 : OAI22_X1 port map( A1 => mult_42_I7_n379, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n380, ZN => mult_42_I7_n114);
   mult_42_I7_U350 : XOR2_X1 port map( A => B(63), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n378);
   mult_42_I7_U349 : OAI22_X1 port map( A1 => mult_42_I7_n378, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n379, ZN => mult_42_I7_n115);
   mult_42_I7_U348 : XOR2_X1 port map( A => B(62), B => mult_42_I7_n314, Z => 
                           mult_42_I7_n377);
   mult_42_I7_U347 : OAI22_X1 port map( A1 => mult_42_I7_n377, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n378, ZN => mult_42_I7_n116);
   mult_42_I7_U346 : XOR2_X1 port map( A => mult_42_I7_n312, B => 
                           x_vector_69_port, Z => mult_42_I7_n376);
   mult_42_I7_U345 : OAI22_X1 port map( A1 => mult_42_I7_n376, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n377, ZN => mult_42_I7_n117);
   mult_42_I7_U344 : XOR2_X1 port map( A => mult_42_I7_n314, B => B(60), Z => 
                           mult_42_I7_n375);
   mult_42_I7_U343 : OAI22_X1 port map( A1 => mult_42_I7_n375, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n376, ZN => mult_42_I7_n118);
   mult_42_I7_U342 : NOR2_X1 port map( A1 => mult_42_I7_n338, A2 => 
                           mult_42_I7_n313, ZN => mult_42_I7_n119);
   mult_42_I7_U341 : XOR2_X1 port map( A => B(69), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n335);
   mult_42_I7_U340 : OAI22_X1 port map( A1 => mult_42_I7_n335, A2 => 
                           mult_42_I7_n327, B1 => mult_42_I7_n326, B2 => 
                           mult_42_I7_n335, ZN => mult_42_I7_n374);
   mult_42_I7_U339 : XOR2_X1 port map( A => B(67), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n373);
   mult_42_I7_U338 : XOR2_X1 port map( A => B(68), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n334);
   mult_42_I7_U337 : OAI22_X1 port map( A1 => mult_42_I7_n373, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n334, ZN => mult_42_I7_n121);
   mult_42_I7_U336 : XOR2_X1 port map( A => B(66), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n372);
   mult_42_I7_U335 : OAI22_X1 port map( A1 => mult_42_I7_n372, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n373, ZN => mult_42_I7_n122);
   mult_42_I7_U334 : XOR2_X1 port map( A => B(65), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n371);
   mult_42_I7_U333 : OAI22_X1 port map( A1 => mult_42_I7_n371, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n372, ZN => mult_42_I7_n123);
   mult_42_I7_U332 : XOR2_X1 port map( A => B(64), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n328);
   mult_42_I7_U331 : OAI22_X1 port map( A1 => mult_42_I7_n328, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n371, ZN => mult_42_I7_n124);
   mult_42_I7_U330 : XOR2_X1 port map( A => B(62), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n370);
   mult_42_I7_U329 : XOR2_X1 port map( A => B(63), B => mult_42_I7_n315, Z => 
                           mult_42_I7_n325);
   mult_42_I7_U328 : OAI22_X1 port map( A1 => mult_42_I7_n370, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n325, ZN => mult_42_I7_n126);
   mult_42_I7_U327 : XOR2_X1 port map( A => mult_42_I7_n312, B => 
                           x_vector_67_port, Z => mult_42_I7_n369);
   mult_42_I7_U326 : OAI22_X1 port map( A1 => mult_42_I7_n369, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n370, ZN => mult_42_I7_n127);
   mult_42_I7_U325 : XOR2_X1 port map( A => mult_42_I7_n313, B => 
                           x_vector_67_port, Z => mult_42_I7_n368);
   mult_42_I7_U324 : OAI22_X1 port map( A1 => mult_42_I7_n368, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n369, ZN => mult_42_I7_n128);
   mult_42_I7_U323 : NOR2_X1 port map( A1 => mult_42_I7_n327, A2 => 
                           mult_42_I7_n313, ZN => mult_42_I7_n129);
   mult_42_I7_U322 : XOR2_X1 port map( A => B(69), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n333);
   mult_42_I7_U321 : OAI22_X1 port map( A1 => mult_42_I7_n333, A2 => 
                           mult_42_I7_n332, B1 => mult_42_I7_n331, B2 => 
                           mult_42_I7_n333, ZN => mult_42_I7_n367);
   mult_42_I7_U320 : XOR2_X1 port map( A => B(67), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n366);
   mult_42_I7_U319 : XOR2_X1 port map( A => B(68), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n330);
   mult_42_I7_U318 : OAI22_X1 port map( A1 => mult_42_I7_n366, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n330, ZN => mult_42_I7_n131);
   mult_42_I7_U317 : XOR2_X1 port map( A => B(66), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n365);
   mult_42_I7_U316 : OAI22_X1 port map( A1 => mult_42_I7_n365, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n366, ZN => mult_42_I7_n132);
   mult_42_I7_U315 : XOR2_X1 port map( A => B(65), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n364);
   mult_42_I7_U314 : OAI22_X1 port map( A1 => mult_42_I7_n364, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n365, ZN => mult_42_I7_n133);
   mult_42_I7_U313 : XOR2_X1 port map( A => B(64), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n363);
   mult_42_I7_U312 : OAI22_X1 port map( A1 => mult_42_I7_n363, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n364, ZN => mult_42_I7_n134);
   mult_42_I7_U311 : XOR2_X1 port map( A => B(63), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n362);
   mult_42_I7_U310 : OAI22_X1 port map( A1 => mult_42_I7_n362, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n363, ZN => mult_42_I7_n135);
   mult_42_I7_U309 : XOR2_X1 port map( A => B(62), B => mult_42_I7_n316, Z => 
                           mult_42_I7_n361);
   mult_42_I7_U308 : OAI22_X1 port map( A1 => mult_42_I7_n361, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n362, ZN => mult_42_I7_n136);
   mult_42_I7_U307 : XOR2_X1 port map( A => mult_42_I7_n312, B => 
                           x_vector_65_port, Z => mult_42_I7_n360);
   mult_42_I7_U306 : OAI22_X1 port map( A1 => mult_42_I7_n360, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n361, ZN => mult_42_I7_n137);
   mult_42_I7_U305 : XOR2_X1 port map( A => mult_42_I7_n313, B => 
                           x_vector_65_port, Z => mult_42_I7_n359);
   mult_42_I7_U304 : OAI22_X1 port map( A1 => mult_42_I7_n359, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n360, ZN => mult_42_I7_n138);
   mult_42_I7_U303 : NOR2_X1 port map( A1 => mult_42_I7_n332, A2 => 
                           mult_42_I7_n313, ZN => mult_42_I7_n139);
   mult_42_I7_U302 : XOR2_X1 port map( A => B(69), B => x_vector_63_port, Z => 
                           mult_42_I7_n329);
   mult_42_I7_U301 : AOI22_X1 port map( A1 => mult_42_I7_n329, A2 => 
                           mult_42_I7_n319, B1 => mult_42_I7_n318, B2 => 
                           mult_42_I7_n329, ZN => mult_42_I7_n140);
   mult_42_I7_U300 : XOR2_X1 port map( A => B(66), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n358);
   mult_42_I7_U299 : XOR2_X1 port map( A => B(67), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n324);
   mult_42_I7_U298 : OAI22_X1 port map( A1 => mult_42_I7_n358, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n324, ZN => mult_42_I7_n142);
   mult_42_I7_U297 : XOR2_X1 port map( A => B(65), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n357);
   mult_42_I7_U296 : OAI22_X1 port map( A1 => mult_42_I7_n357, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n358, ZN => mult_42_I7_n143);
   mult_42_I7_U295 : XOR2_X1 port map( A => B(64), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n356);
   mult_42_I7_U294 : OAI22_X1 port map( A1 => mult_42_I7_n356, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n357, ZN => mult_42_I7_n144);
   mult_42_I7_U293 : XOR2_X1 port map( A => B(63), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n355);
   mult_42_I7_U292 : OAI22_X1 port map( A1 => mult_42_I7_n355, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n356, ZN => mult_42_I7_n145);
   mult_42_I7_U291 : XOR2_X1 port map( A => B(62), B => mult_42_I7_n317, Z => 
                           mult_42_I7_n354);
   mult_42_I7_U290 : OAI22_X1 port map( A1 => mult_42_I7_n354, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n355, ZN => mult_42_I7_n146);
   mult_42_I7_U289 : XOR2_X1 port map( A => mult_42_I7_n312, B => 
                           x_vector_63_port, Z => mult_42_I7_n353);
   mult_42_I7_U288 : OAI22_X1 port map( A1 => mult_42_I7_n353, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n354, ZN => mult_42_I7_n147);
   mult_42_I7_U287 : XOR2_X1 port map( A => mult_42_I7_n313, B => 
                           x_vector_63_port, Z => mult_42_I7_n350);
   mult_42_I7_U286 : OAI22_X1 port map( A1 => mult_42_I7_n350, A2 => 
                           mult_42_I7_n351, B1 => mult_42_I7_n352, B2 => 
                           mult_42_I7_n353, ZN => mult_42_I7_n148);
   mult_42_I7_U285 : XNOR2_X1 port map( A => B(69), B => x_vector_61_port, ZN 
                           => mult_42_I7_n348);
   mult_42_I7_U284 : OAI22_X1 port map( A1 => mult_42_I7_n320, A2 => 
                           mult_42_I7_n348, B1 => mult_42_I7_n341, B2 => 
                           mult_42_I7_n348, ZN => mult_42_I7_n349);
   mult_42_I7_U283 : XNOR2_X1 port map( A => B(68), B => x_vector_61_port, ZN 
                           => mult_42_I7_n347);
   mult_42_I7_U282 : OAI22_X1 port map( A1 => mult_42_I7_n347, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n348, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n151);
   mult_42_I7_U281 : XNOR2_X1 port map( A => B(67), B => x_vector_61_port, ZN 
                           => mult_42_I7_n346);
   mult_42_I7_U280 : OAI22_X1 port map( A1 => mult_42_I7_n346, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n347, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n152);
   mult_42_I7_U279 : XNOR2_X1 port map( A => B(66), B => x_vector_61_port, ZN 
                           => mult_42_I7_n345);
   mult_42_I7_U278 : OAI22_X1 port map( A1 => mult_42_I7_n345, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n346, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n153);
   mult_42_I7_U277 : XNOR2_X1 port map( A => B(65), B => x_vector_61_port, ZN 
                           => mult_42_I7_n344);
   mult_42_I7_U276 : OAI22_X1 port map( A1 => mult_42_I7_n344, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n345, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n154);
   mult_42_I7_U275 : XNOR2_X1 port map( A => B(64), B => x_vector_61_port, ZN 
                           => mult_42_I7_n343);
   mult_42_I7_U274 : OAI22_X1 port map( A1 => mult_42_I7_n343, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n344, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n155);
   mult_42_I7_U273 : XNOR2_X1 port map( A => B(63), B => x_vector_61_port, ZN 
                           => mult_42_I7_n342);
   mult_42_I7_U272 : OAI22_X1 port map( A1 => mult_42_I7_n342, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n343, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n156);
   mult_42_I7_U271 : OAI22_X1 port map( A1 => mult_42_I7_n340, A2 => 
                           mult_42_I7_n341, B1 => mult_42_I7_n342, B2 => 
                           mult_42_I7_n320, ZN => mult_42_I7_n157);
   mult_42_I7_U270 : OAI22_X1 port map( A1 => mult_42_I7_n336, A2 => 
                           mult_42_I7_n337, B1 => mult_42_I7_n338, B2 => 
                           mult_42_I7_n339, ZN => mult_42_I7_n19);
   mult_42_I7_U269 : OAI22_X1 port map( A1 => mult_42_I7_n334, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n335, ZN => mult_42_I7_n25);
   mult_42_I7_U268 : OAI22_X1 port map( A1 => mult_42_I7_n330, A2 => 
                           mult_42_I7_n331, B1 => mult_42_I7_n332, B2 => 
                           mult_42_I7_n333, ZN => mult_42_I7_n35);
   mult_42_I7_U267 : XOR2_X1 port map( A => B(68), B => x_vector_63_port, Z => 
                           mult_42_I7_n323);
   mult_42_I7_U266 : AOI22_X1 port map( A1 => mult_42_I7_n323, A2 => 
                           mult_42_I7_n318, B1 => mult_42_I7_n319, B2 => 
                           mult_42_I7_n329, ZN => mult_42_I7_n50);
   mult_42_I7_U265 : OAI22_X1 port map( A1 => mult_42_I7_n325, A2 => 
                           mult_42_I7_n326, B1 => mult_42_I7_n327, B2 => 
                           mult_42_I7_n328, ZN => mult_42_I7_n321);
   mult_42_I7_U264 : AOI22_X1 port map( A1 => mult_42_I7_n306, A2 => 
                           mult_42_I7_n318, B1 => mult_42_I7_n319, B2 => 
                           mult_42_I7_n323, ZN => mult_42_I7_n322);
   mult_42_I7_U263 : NAND2_X1 port map( A1 => mult_42_I7_n310, A2 => 
                           mult_42_I7_n322, ZN => mult_42_I7_n57);
   mult_42_I7_U262 : XOR2_X1 port map( A => mult_42_I7_n321, B => 
                           mult_42_I7_n322, Z => mult_42_I7_n58);
   mult_42_I7_U261 : XNOR2_X2 port map( A => x_vector_68_port, B => 
                           x_vector_67_port, ZN => mult_42_I7_n338);
   mult_42_I7_U260 : XNOR2_X2 port map( A => x_vector_66_port, B => 
                           x_vector_65_port, ZN => mult_42_I7_n327);
   mult_42_I7_U259 : XNOR2_X2 port map( A => x_vector_64_port, B => 
                           x_vector_63_port, ZN => mult_42_I7_n332);
   mult_42_I7_U258 : INV_X1 port map( A => B(61), ZN => mult_42_I7_n312);
   mult_42_I7_U257 : INV_X1 port map( A => B(60), ZN => mult_42_I7_n313);
   mult_42_I7_U256 : INV_X1 port map( A => x_vector_63_port, ZN => 
                           mult_42_I7_n317);
   mult_42_I7_U255 : INV_X1 port map( A => x_vector_60_port, ZN => 
                           mult_42_I7_n320);
   mult_42_I7_U254 : INV_X1 port map( A => x_vector_67_port, ZN => 
                           mult_42_I7_n315);
   mult_42_I7_U253 : INV_X1 port map( A => x_vector_65_port, ZN => 
                           mult_42_I7_n316);
   mult_42_I7_U252 : INV_X1 port map( A => x_vector_69_port, ZN => 
                           mult_42_I7_n314);
   mult_42_I7_U251 : INV_X1 port map( A => mult_42_I7_n374, ZN => 
                           mult_42_I7_n300);
   mult_42_I7_U250 : INV_X1 port map( A => mult_42_I7_n25, ZN => 
                           mult_42_I7_n301);
   mult_42_I7_U249 : INV_X1 port map( A => mult_42_I7_n90, ZN => 
                           mult_42_I7_n311);
   mult_42_I7_U248 : INV_X1 port map( A => mult_42_I7_n50, ZN => 
                           mult_42_I7_n297);
   mult_42_I7_U247 : INV_X1 port map( A => mult_42_I7_n367, ZN => 
                           mult_42_I7_n298);
   mult_42_I7_U246 : INV_X1 port map( A => mult_42_I7_n383, ZN => 
                           mult_42_I7_n302);
   mult_42_I7_U245 : INV_X1 port map( A => mult_42_I7_n349, ZN => 
                           mult_42_I7_n295);
   mult_42_I7_U244 : INV_X1 port map( A => mult_42_I7_n35, ZN => 
                           mult_42_I7_n299);
   mult_42_I7_U243 : INV_X1 port map( A => mult_42_I7_n351, ZN => 
                           mult_42_I7_n318);
   mult_42_I7_U242 : INV_X1 port map( A => mult_42_I7_n352, ZN => 
                           mult_42_I7_n319);
   mult_42_I7_U241 : INV_X1 port map( A => mult_42_I7_n324, ZN => 
                           mult_42_I7_n306);
   mult_42_I7_U240 : INV_X1 port map( A => mult_42_I7_n84, ZN => 
                           mult_42_I7_n308);
   mult_42_I7_U239 : INV_X1 port map( A => mult_42_I7_n87, ZN => 
                           mult_42_I7_n309);
   mult_42_I7_U238 : INV_X1 port map( A => mult_42_I7_n19, ZN => 
                           mult_42_I7_n303);
   mult_42_I7_U237 : INV_X1 port map( A => mult_42_I7_n321, ZN => 
                           mult_42_I7_n310);
   mult_42_I7_U236 : INV_X1 port map( A => mult_42_I7_n1, ZN => N122);
   mult_42_I7_U235 : INV_X1 port map( A => mult_42_I7_n74, ZN => 
                           mult_42_I7_n305);
   mult_42_I7_U234 : INV_X1 port map( A => mult_42_I7_n79, ZN => 
                           mult_42_I7_n307);
   mult_42_I7_U233 : INV_X1 port map( A => mult_42_I7_n60, ZN => 
                           mult_42_I7_n296);
   mult_42_I7_U232 : INV_X1 port map( A => mult_42_I7_n67, ZN => 
                           mult_42_I7_n304);
   mult_42_I7_U56 : HA_X1 port map( A => mult_42_I7_n148, B => mult_42_I7_n157,
                           CO => mult_42_I7_n89, S => mult_42_I7_n90);
   mult_42_I7_U55 : FA_X1 port map( A => mult_42_I7_n156, B => mult_42_I7_n139,
                           CI => mult_42_I7_n147, CO => mult_42_I7_n87, S => 
                           mult_42_I7_n88);
   mult_42_I7_U54 : HA_X1 port map( A => mult_42_I7_n107, B => mult_42_I7_n138,
                           CO => mult_42_I7_n85, S => mult_42_I7_n86);
   mult_42_I7_U53 : FA_X1 port map( A => mult_42_I7_n146, B => mult_42_I7_n155,
                           CI => mult_42_I7_n86, CO => mult_42_I7_n83, S => 
                           mult_42_I7_n84);
   mult_42_I7_U52 : FA_X1 port map( A => mult_42_I7_n154, B => mult_42_I7_n129,
                           CI => mult_42_I7_n145, CO => mult_42_I7_n81, S => 
                           mult_42_I7_n82);
   mult_42_I7_U51 : FA_X1 port map( A => mult_42_I7_n85, B => mult_42_I7_n137, 
                           CI => mult_42_I7_n82, CO => mult_42_I7_n79, S => 
                           mult_42_I7_n80);
   mult_42_I7_U50 : HA_X1 port map( A => mult_42_I7_n106, B => mult_42_I7_n128,
                           CO => mult_42_I7_n77, S => mult_42_I7_n78);
   mult_42_I7_U49 : FA_X1 port map( A => mult_42_I7_n136, B => mult_42_I7_n153,
                           CI => mult_42_I7_n144, CO => mult_42_I7_n75, S => 
                           mult_42_I7_n76);
   mult_42_I7_U48 : FA_X1 port map( A => mult_42_I7_n81, B => mult_42_I7_n78, 
                           CI => mult_42_I7_n76, CO => mult_42_I7_n73, S => 
                           mult_42_I7_n74);
   mult_42_I7_U47 : FA_X1 port map( A => mult_42_I7_n135, B => mult_42_I7_n119,
                           CI => mult_42_I7_n152, CO => mult_42_I7_n71, S => 
                           mult_42_I7_n72);
   mult_42_I7_U46 : FA_X1 port map( A => mult_42_I7_n127, B => mult_42_I7_n143,
                           CI => mult_42_I7_n77, CO => mult_42_I7_n69, S => 
                           mult_42_I7_n70);
   mult_42_I7_U45 : FA_X1 port map( A => mult_42_I7_n72, B => mult_42_I7_n75, 
                           CI => mult_42_I7_n70, CO => mult_42_I7_n67, S => 
                           mult_42_I7_n68);
   mult_42_I7_U44 : HA_X1 port map( A => mult_42_I7_n105, B => mult_42_I7_n118,
                           CO => mult_42_I7_n65, S => mult_42_I7_n66);
   mult_42_I7_U43 : FA_X1 port map( A => mult_42_I7_n126, B => mult_42_I7_n134,
                           CI => mult_42_I7_n142, CO => mult_42_I7_n63, S => 
                           mult_42_I7_n64);
   mult_42_I7_U42 : FA_X1 port map( A => mult_42_I7_n66, B => mult_42_I7_n151, 
                           CI => mult_42_I7_n71, CO => mult_42_I7_n61, S => 
                           mult_42_I7_n62);
   mult_42_I7_U41 : FA_X1 port map( A => mult_42_I7_n64, B => mult_42_I7_n69, 
                           CI => mult_42_I7_n62, CO => mult_42_I7_n59, S => 
                           mult_42_I7_n60);
   mult_42_I7_U38 : FA_X1 port map( A => mult_42_I7_n133, B => mult_42_I7_n117,
                           CI => mult_42_I7_n295, CO => mult_42_I7_n55, S => 
                           mult_42_I7_n56);
   mult_42_I7_U37 : FA_X1 port map( A => mult_42_I7_n58, B => mult_42_I7_n65, 
                           CI => mult_42_I7_n63, CO => mult_42_I7_n53, S => 
                           mult_42_I7_n54);
   mult_42_I7_U36 : FA_X1 port map( A => mult_42_I7_n61, B => mult_42_I7_n56, 
                           CI => mult_42_I7_n54, CO => mult_42_I7_n51, S => 
                           mult_42_I7_n52);
   mult_42_I7_U34 : FA_X1 port map( A => mult_42_I7_n124, B => mult_42_I7_n116,
                           CI => mult_42_I7_n132, CO => mult_42_I7_n47, S => 
                           mult_42_I7_n48);
   mult_42_I7_U33 : FA_X1 port map( A => mult_42_I7_n57, B => mult_42_I7_n50, 
                           CI => mult_42_I7_n55, CO => mult_42_I7_n45, S => 
                           mult_42_I7_n46);
   mult_42_I7_U32 : FA_X1 port map( A => mult_42_I7_n53, B => mult_42_I7_n48, 
                           CI => mult_42_I7_n46, CO => mult_42_I7_n43, S => 
                           mult_42_I7_n44);
   mult_42_I7_U31 : FA_X1 port map( A => mult_42_I7_n123, B => mult_42_I7_n115,
                           CI => mult_42_I7_n140, CO => mult_42_I7_n41, S => 
                           mult_42_I7_n42);
   mult_42_I7_U30 : FA_X1 port map( A => mult_42_I7_n297, B => mult_42_I7_n131,
                           CI => mult_42_I7_n47, CO => mult_42_I7_n39, S => 
                           mult_42_I7_n40);
   mult_42_I7_U29 : FA_X1 port map( A => mult_42_I7_n45, B => mult_42_I7_n42, 
                           CI => mult_42_I7_n40, CO => mult_42_I7_n37, S => 
                           mult_42_I7_n38);
   mult_42_I7_U27 : FA_X1 port map( A => mult_42_I7_n114, B => mult_42_I7_n122,
                           CI => mult_42_I7_n299, CO => mult_42_I7_n33, S => 
                           mult_42_I7_n34);
   mult_42_I7_U26 : FA_X1 port map( A => mult_42_I7_n34, B => mult_42_I7_n41, 
                           CI => mult_42_I7_n39, CO => mult_42_I7_n31, S => 
                           mult_42_I7_n32);
   mult_42_I7_U25 : FA_X1 port map( A => mult_42_I7_n121, B => mult_42_I7_n35, 
                           CI => mult_42_I7_n298, CO => mult_42_I7_n29, S => 
                           mult_42_I7_n30);
   mult_42_I7_U24 : FA_X1 port map( A => mult_42_I7_n33, B => mult_42_I7_n113, 
                           CI => mult_42_I7_n30, CO => mult_42_I7_n27, S => 
                           mult_42_I7_n28);
   mult_42_I7_U22 : FA_X1 port map( A => mult_42_I7_n301, B => mult_42_I7_n112,
                           CI => mult_42_I7_n29, CO => mult_42_I7_n23, S => 
                           mult_42_I7_n24);
   mult_42_I7_U21 : FA_X1 port map( A => mult_42_I7_n111, B => mult_42_I7_n25, 
                           CI => mult_42_I7_n300, CO => mult_42_I7_n21, S => 
                           mult_42_I7_n22);
   mult_42_I7_U10 : FA_X1 port map( A => mult_42_I7_n52, B => mult_42_I7_n59, 
                           CI => mult_42_I7_n10, CO => mult_42_I7_n9, S => N113
                           );
   mult_42_I7_U9 : FA_X1 port map( A => mult_42_I7_n44, B => mult_42_I7_n51, CI
                           => mult_42_I7_n9, CO => mult_42_I7_n8, S => N114);
   mult_42_I7_U8 : FA_X1 port map( A => mult_42_I7_n38, B => mult_42_I7_n43, CI
                           => mult_42_I7_n8, CO => mult_42_I7_n7, S => N115);
   mult_42_I7_U7 : FA_X1 port map( A => mult_42_I7_n32, B => mult_42_I7_n37, CI
                           => mult_42_I7_n7, CO => mult_42_I7_n6, S => N116);
   mult_42_I7_U6 : FA_X1 port map( A => mult_42_I7_n28, B => mult_42_I7_n31, CI
                           => mult_42_I7_n6, CO => mult_42_I7_n5, S => N117);
   mult_42_I7_U5 : FA_X1 port map( A => mult_42_I7_n24, B => mult_42_I7_n27, CI
                           => mult_42_I7_n5, CO => mult_42_I7_n4, S => N118);
   mult_42_I7_U4 : FA_X1 port map( A => mult_42_I7_n23, B => mult_42_I7_n22, CI
                           => mult_42_I7_n4, CO => mult_42_I7_n3, S => N119);
   mult_42_I7_U3 : FA_X1 port map( A => mult_42_I7_n21, B => mult_42_I7_n303, 
                           CI => mult_42_I7_n3, CO => mult_42_I7_n2, S => N120)
                           ;
   mult_42_I7_U2 : FA_X1 port map( A => mult_42_I7_n302, B => mult_42_I7_n19, 
                           CI => mult_42_I7_n2, CO => mult_42_I7_n1, S => N121)
                           ;
   mult_42_I8_U391 : NAND2_X1 port map( A1 => x_vector_71_port, A2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n341);
   mult_42_I8_U390 : XNOR2_X1 port map( A => B(72), B => x_vector_71_port, ZN 
                           => mult_42_I8_n340);
   mult_42_I8_U389 : OAI22_X1 port map( A1 => B(71), A2 => mult_42_I8_n341, B1 
                           => mult_42_I8_n340, B2 => mult_42_I8_n320, ZN => 
                           mult_42_I8_n402);
   mult_42_I8_U388 : NAND3_X1 port map( A1 => mult_42_I8_n402, A2 => 
                           mult_42_I8_n312, A3 => x_vector_71_port, ZN => 
                           mult_42_I8_n400);
   mult_42_I8_U387 : XNOR2_X1 port map( A => x_vector_72_port, B => 
                           x_vector_71_port, ZN => mult_42_I8_n352);
   mult_42_I8_U386 : NAND2_X1 port map( A1 => mult_42_I8_n319, A2 => 
                           mult_42_I8_n402, ZN => mult_42_I8_n401);
   mult_42_I8_U385 : MUX2_X1 port map( A => mult_42_I8_n400, B => 
                           mult_42_I8_n401, S => B(70), Z => mult_42_I8_n396);
   mult_42_I8_U384 : XOR2_X1 port map( A => x_vector_73_port, B => 
                           x_vector_72_port, Z => mult_42_I8_n399);
   mult_42_I8_U383 : NAND2_X1 port map( A1 => mult_42_I8_n352, A2 => 
                           mult_42_I8_n399, ZN => mult_42_I8_n351);
   mult_42_I8_U382 : NOR3_X1 port map( A1 => mult_42_I8_n352, A2 => B(70), A3 
                           => mult_42_I8_n317, ZN => mult_42_I8_n398);
   mult_42_I8_U381 : AOI21_X1 port map( B1 => x_vector_73_port, B2 => 
                           mult_42_I8_n318, A => mult_42_I8_n398, ZN => 
                           mult_42_I8_n397);
   mult_42_I8_U380 : OAI222_X1 port map( A1 => mult_42_I8_n396, A2 => 
                           mult_42_I8_n311, B1 => mult_42_I8_n397, B2 => 
                           mult_42_I8_n396, C1 => mult_42_I8_n397, C2 => 
                           mult_42_I8_n311, ZN => mult_42_I8_n395);
   mult_42_I8_U379 : AOI222_X1 port map( A1 => mult_42_I8_n395, A2 => 
                           mult_42_I8_n88, B1 => mult_42_I8_n395, B2 => 
                           mult_42_I8_n89, C1 => mult_42_I8_n89, C2 => 
                           mult_42_I8_n88, ZN => mult_42_I8_n394);
   mult_42_I8_U378 : OAI222_X1 port map( A1 => mult_42_I8_n394, A2 => 
                           mult_42_I8_n308, B1 => mult_42_I8_n394, B2 => 
                           mult_42_I8_n309, C1 => mult_42_I8_n309, C2 => 
                           mult_42_I8_n308, ZN => mult_42_I8_n393);
   mult_42_I8_U377 : AOI222_X1 port map( A1 => mult_42_I8_n393, A2 => 
                           mult_42_I8_n80, B1 => mult_42_I8_n393, B2 => 
                           mult_42_I8_n83, C1 => mult_42_I8_n83, C2 => 
                           mult_42_I8_n80, ZN => mult_42_I8_n392);
   mult_42_I8_U376 : OAI222_X1 port map( A1 => mult_42_I8_n392, A2 => 
                           mult_42_I8_n305, B1 => mult_42_I8_n392, B2 => 
                           mult_42_I8_n307, C1 => mult_42_I8_n307, C2 => 
                           mult_42_I8_n305, ZN => mult_42_I8_n391);
   mult_42_I8_U375 : AOI222_X1 port map( A1 => mult_42_I8_n391, A2 => 
                           mult_42_I8_n68, B1 => mult_42_I8_n391, B2 => 
                           mult_42_I8_n73, C1 => mult_42_I8_n73, C2 => 
                           mult_42_I8_n68, ZN => mult_42_I8_n390);
   mult_42_I8_U374 : OAI222_X1 port map( A1 => mult_42_I8_n390, A2 => 
                           mult_42_I8_n296, B1 => mult_42_I8_n390, B2 => 
                           mult_42_I8_n304, C1 => mult_42_I8_n304, C2 => 
                           mult_42_I8_n296, ZN => mult_42_I8_n10);
   mult_42_I8_U373 : XOR2_X1 port map( A => x_vector_79_port, B => 
                           x_vector_78_port, Z => mult_42_I8_n389);
   mult_42_I8_U372 : NAND2_X1 port map( A1 => mult_42_I8_n338, A2 => 
                           mult_42_I8_n389, ZN => mult_42_I8_n337);
   mult_42_I8_U371 : OR3_X1 port map( A1 => mult_42_I8_n338, A2 => B(70), A3 =>
                           mult_42_I8_n314, ZN => mult_42_I8_n388);
   mult_42_I8_U370 : OAI21_X1 port map( B1 => mult_42_I8_n314, B2 => 
                           mult_42_I8_n337, A => mult_42_I8_n388, ZN => 
                           mult_42_I8_n105);
   mult_42_I8_U369 : XOR2_X1 port map( A => x_vector_77_port, B => 
                           x_vector_76_port, Z => mult_42_I8_n387);
   mult_42_I8_U368 : NAND2_X1 port map( A1 => mult_42_I8_n327, A2 => 
                           mult_42_I8_n387, ZN => mult_42_I8_n326);
   mult_42_I8_U367 : OR3_X1 port map( A1 => mult_42_I8_n327, A2 => B(70), A3 =>
                           mult_42_I8_n315, ZN => mult_42_I8_n386);
   mult_42_I8_U366 : OAI21_X1 port map( B1 => mult_42_I8_n315, B2 => 
                           mult_42_I8_n326, A => mult_42_I8_n386, ZN => 
                           mult_42_I8_n106);
   mult_42_I8_U365 : XOR2_X1 port map( A => x_vector_75_port, B => 
                           x_vector_74_port, Z => mult_42_I8_n385);
   mult_42_I8_U364 : NAND2_X1 port map( A1 => mult_42_I8_n332, A2 => 
                           mult_42_I8_n385, ZN => mult_42_I8_n331);
   mult_42_I8_U363 : OR3_X1 port map( A1 => mult_42_I8_n332, A2 => B(70), A3 =>
                           mult_42_I8_n316, ZN => mult_42_I8_n384);
   mult_42_I8_U362 : OAI21_X1 port map( B1 => mult_42_I8_n316, B2 => 
                           mult_42_I8_n331, A => mult_42_I8_n384, ZN => 
                           mult_42_I8_n107);
   mult_42_I8_U361 : XOR2_X1 port map( A => B(79), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n339);
   mult_42_I8_U360 : OAI22_X1 port map( A1 => mult_42_I8_n339, A2 => 
                           mult_42_I8_n338, B1 => mult_42_I8_n337, B2 => 
                           mult_42_I8_n339, ZN => mult_42_I8_n383);
   mult_42_I8_U359 : XOR2_X1 port map( A => B(77), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n382);
   mult_42_I8_U358 : XOR2_X1 port map( A => B(78), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n336);
   mult_42_I8_U357 : OAI22_X1 port map( A1 => mult_42_I8_n382, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n336, ZN => mult_42_I8_n111);
   mult_42_I8_U356 : XOR2_X1 port map( A => B(76), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n381);
   mult_42_I8_U355 : OAI22_X1 port map( A1 => mult_42_I8_n381, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n382, ZN => mult_42_I8_n112);
   mult_42_I8_U354 : XOR2_X1 port map( A => B(75), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n380);
   mult_42_I8_U353 : OAI22_X1 port map( A1 => mult_42_I8_n380, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n381, ZN => mult_42_I8_n113);
   mult_42_I8_U352 : XOR2_X1 port map( A => B(74), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n379);
   mult_42_I8_U351 : OAI22_X1 port map( A1 => mult_42_I8_n379, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n380, ZN => mult_42_I8_n114);
   mult_42_I8_U350 : XOR2_X1 port map( A => B(73), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n378);
   mult_42_I8_U349 : OAI22_X1 port map( A1 => mult_42_I8_n378, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n379, ZN => mult_42_I8_n115);
   mult_42_I8_U348 : XOR2_X1 port map( A => B(72), B => mult_42_I8_n314, Z => 
                           mult_42_I8_n377);
   mult_42_I8_U347 : OAI22_X1 port map( A1 => mult_42_I8_n377, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n378, ZN => mult_42_I8_n116);
   mult_42_I8_U346 : XOR2_X1 port map( A => mult_42_I8_n312, B => 
                           x_vector_79_port, Z => mult_42_I8_n376);
   mult_42_I8_U345 : OAI22_X1 port map( A1 => mult_42_I8_n376, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n377, ZN => mult_42_I8_n117);
   mult_42_I8_U344 : XOR2_X1 port map( A => mult_42_I8_n314, B => B(70), Z => 
                           mult_42_I8_n375);
   mult_42_I8_U343 : OAI22_X1 port map( A1 => mult_42_I8_n375, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n376, ZN => mult_42_I8_n118);
   mult_42_I8_U342 : NOR2_X1 port map( A1 => mult_42_I8_n338, A2 => 
                           mult_42_I8_n313, ZN => mult_42_I8_n119);
   mult_42_I8_U341 : XOR2_X1 port map( A => B(79), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n335);
   mult_42_I8_U340 : OAI22_X1 port map( A1 => mult_42_I8_n335, A2 => 
                           mult_42_I8_n327, B1 => mult_42_I8_n326, B2 => 
                           mult_42_I8_n335, ZN => mult_42_I8_n374);
   mult_42_I8_U339 : XOR2_X1 port map( A => B(77), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n373);
   mult_42_I8_U338 : XOR2_X1 port map( A => B(78), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n334);
   mult_42_I8_U337 : OAI22_X1 port map( A1 => mult_42_I8_n373, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n334, ZN => mult_42_I8_n121);
   mult_42_I8_U336 : XOR2_X1 port map( A => B(76), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n372);
   mult_42_I8_U335 : OAI22_X1 port map( A1 => mult_42_I8_n372, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n373, ZN => mult_42_I8_n122);
   mult_42_I8_U334 : XOR2_X1 port map( A => B(75), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n371);
   mult_42_I8_U333 : OAI22_X1 port map( A1 => mult_42_I8_n371, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n372, ZN => mult_42_I8_n123);
   mult_42_I8_U332 : XOR2_X1 port map( A => B(74), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n328);
   mult_42_I8_U331 : OAI22_X1 port map( A1 => mult_42_I8_n328, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n371, ZN => mult_42_I8_n124);
   mult_42_I8_U330 : XOR2_X1 port map( A => B(72), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n370);
   mult_42_I8_U329 : XOR2_X1 port map( A => B(73), B => mult_42_I8_n315, Z => 
                           mult_42_I8_n325);
   mult_42_I8_U328 : OAI22_X1 port map( A1 => mult_42_I8_n370, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n325, ZN => mult_42_I8_n126);
   mult_42_I8_U327 : XOR2_X1 port map( A => mult_42_I8_n312, B => 
                           x_vector_77_port, Z => mult_42_I8_n369);
   mult_42_I8_U326 : OAI22_X1 port map( A1 => mult_42_I8_n369, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n370, ZN => mult_42_I8_n127);
   mult_42_I8_U325 : XOR2_X1 port map( A => mult_42_I8_n313, B => 
                           x_vector_77_port, Z => mult_42_I8_n368);
   mult_42_I8_U324 : OAI22_X1 port map( A1 => mult_42_I8_n368, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n369, ZN => mult_42_I8_n128);
   mult_42_I8_U323 : NOR2_X1 port map( A1 => mult_42_I8_n327, A2 => 
                           mult_42_I8_n313, ZN => mult_42_I8_n129);
   mult_42_I8_U322 : XOR2_X1 port map( A => B(79), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n333);
   mult_42_I8_U321 : OAI22_X1 port map( A1 => mult_42_I8_n333, A2 => 
                           mult_42_I8_n332, B1 => mult_42_I8_n331, B2 => 
                           mult_42_I8_n333, ZN => mult_42_I8_n367);
   mult_42_I8_U320 : XOR2_X1 port map( A => B(77), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n366);
   mult_42_I8_U319 : XOR2_X1 port map( A => B(78), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n330);
   mult_42_I8_U318 : OAI22_X1 port map( A1 => mult_42_I8_n366, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n330, ZN => mult_42_I8_n131);
   mult_42_I8_U317 : XOR2_X1 port map( A => B(76), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n365);
   mult_42_I8_U316 : OAI22_X1 port map( A1 => mult_42_I8_n365, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n366, ZN => mult_42_I8_n132);
   mult_42_I8_U315 : XOR2_X1 port map( A => B(75), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n364);
   mult_42_I8_U314 : OAI22_X1 port map( A1 => mult_42_I8_n364, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n365, ZN => mult_42_I8_n133);
   mult_42_I8_U313 : XOR2_X1 port map( A => B(74), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n363);
   mult_42_I8_U312 : OAI22_X1 port map( A1 => mult_42_I8_n363, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n364, ZN => mult_42_I8_n134);
   mult_42_I8_U311 : XOR2_X1 port map( A => B(73), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n362);
   mult_42_I8_U310 : OAI22_X1 port map( A1 => mult_42_I8_n362, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n363, ZN => mult_42_I8_n135);
   mult_42_I8_U309 : XOR2_X1 port map( A => B(72), B => mult_42_I8_n316, Z => 
                           mult_42_I8_n361);
   mult_42_I8_U308 : OAI22_X1 port map( A1 => mult_42_I8_n361, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n362, ZN => mult_42_I8_n136);
   mult_42_I8_U307 : XOR2_X1 port map( A => mult_42_I8_n312, B => 
                           x_vector_75_port, Z => mult_42_I8_n360);
   mult_42_I8_U306 : OAI22_X1 port map( A1 => mult_42_I8_n360, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n361, ZN => mult_42_I8_n137);
   mult_42_I8_U305 : XOR2_X1 port map( A => mult_42_I8_n313, B => 
                           x_vector_75_port, Z => mult_42_I8_n359);
   mult_42_I8_U304 : OAI22_X1 port map( A1 => mult_42_I8_n359, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n360, ZN => mult_42_I8_n138);
   mult_42_I8_U303 : NOR2_X1 port map( A1 => mult_42_I8_n332, A2 => 
                           mult_42_I8_n313, ZN => mult_42_I8_n139);
   mult_42_I8_U302 : XOR2_X1 port map( A => B(79), B => x_vector_73_port, Z => 
                           mult_42_I8_n329);
   mult_42_I8_U301 : AOI22_X1 port map( A1 => mult_42_I8_n329, A2 => 
                           mult_42_I8_n319, B1 => mult_42_I8_n318, B2 => 
                           mult_42_I8_n329, ZN => mult_42_I8_n140);
   mult_42_I8_U300 : XOR2_X1 port map( A => B(76), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n358);
   mult_42_I8_U299 : XOR2_X1 port map( A => B(77), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n324);
   mult_42_I8_U298 : OAI22_X1 port map( A1 => mult_42_I8_n358, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n324, ZN => mult_42_I8_n142);
   mult_42_I8_U297 : XOR2_X1 port map( A => B(75), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n357);
   mult_42_I8_U296 : OAI22_X1 port map( A1 => mult_42_I8_n357, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n358, ZN => mult_42_I8_n143);
   mult_42_I8_U295 : XOR2_X1 port map( A => B(74), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n356);
   mult_42_I8_U294 : OAI22_X1 port map( A1 => mult_42_I8_n356, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n357, ZN => mult_42_I8_n144);
   mult_42_I8_U293 : XOR2_X1 port map( A => B(73), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n355);
   mult_42_I8_U292 : OAI22_X1 port map( A1 => mult_42_I8_n355, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n356, ZN => mult_42_I8_n145);
   mult_42_I8_U291 : XOR2_X1 port map( A => B(72), B => mult_42_I8_n317, Z => 
                           mult_42_I8_n354);
   mult_42_I8_U290 : OAI22_X1 port map( A1 => mult_42_I8_n354, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n355, ZN => mult_42_I8_n146);
   mult_42_I8_U289 : XOR2_X1 port map( A => mult_42_I8_n312, B => 
                           x_vector_73_port, Z => mult_42_I8_n353);
   mult_42_I8_U288 : OAI22_X1 port map( A1 => mult_42_I8_n353, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n354, ZN => mult_42_I8_n147);
   mult_42_I8_U287 : XOR2_X1 port map( A => mult_42_I8_n313, B => 
                           x_vector_73_port, Z => mult_42_I8_n350);
   mult_42_I8_U286 : OAI22_X1 port map( A1 => mult_42_I8_n350, A2 => 
                           mult_42_I8_n351, B1 => mult_42_I8_n352, B2 => 
                           mult_42_I8_n353, ZN => mult_42_I8_n148);
   mult_42_I8_U285 : XNOR2_X1 port map( A => B(79), B => x_vector_71_port, ZN 
                           => mult_42_I8_n348);
   mult_42_I8_U284 : OAI22_X1 port map( A1 => mult_42_I8_n320, A2 => 
                           mult_42_I8_n348, B1 => mult_42_I8_n341, B2 => 
                           mult_42_I8_n348, ZN => mult_42_I8_n349);
   mult_42_I8_U283 : XNOR2_X1 port map( A => B(78), B => x_vector_71_port, ZN 
                           => mult_42_I8_n347);
   mult_42_I8_U282 : OAI22_X1 port map( A1 => mult_42_I8_n347, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n348, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n151);
   mult_42_I8_U281 : XNOR2_X1 port map( A => B(77), B => x_vector_71_port, ZN 
                           => mult_42_I8_n346);
   mult_42_I8_U280 : OAI22_X1 port map( A1 => mult_42_I8_n346, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n347, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n152);
   mult_42_I8_U279 : XNOR2_X1 port map( A => B(76), B => x_vector_71_port, ZN 
                           => mult_42_I8_n345);
   mult_42_I8_U278 : OAI22_X1 port map( A1 => mult_42_I8_n345, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n346, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n153);
   mult_42_I8_U277 : XNOR2_X1 port map( A => B(75), B => x_vector_71_port, ZN 
                           => mult_42_I8_n344);
   mult_42_I8_U276 : OAI22_X1 port map( A1 => mult_42_I8_n344, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n345, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n154);
   mult_42_I8_U275 : XNOR2_X1 port map( A => B(74), B => x_vector_71_port, ZN 
                           => mult_42_I8_n343);
   mult_42_I8_U274 : OAI22_X1 port map( A1 => mult_42_I8_n343, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n344, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n155);
   mult_42_I8_U273 : XNOR2_X1 port map( A => B(73), B => x_vector_71_port, ZN 
                           => mult_42_I8_n342);
   mult_42_I8_U272 : OAI22_X1 port map( A1 => mult_42_I8_n342, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n343, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n156);
   mult_42_I8_U271 : OAI22_X1 port map( A1 => mult_42_I8_n340, A2 => 
                           mult_42_I8_n341, B1 => mult_42_I8_n342, B2 => 
                           mult_42_I8_n320, ZN => mult_42_I8_n157);
   mult_42_I8_U270 : OAI22_X1 port map( A1 => mult_42_I8_n336, A2 => 
                           mult_42_I8_n337, B1 => mult_42_I8_n338, B2 => 
                           mult_42_I8_n339, ZN => mult_42_I8_n19);
   mult_42_I8_U269 : OAI22_X1 port map( A1 => mult_42_I8_n334, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n335, ZN => mult_42_I8_n25);
   mult_42_I8_U268 : OAI22_X1 port map( A1 => mult_42_I8_n330, A2 => 
                           mult_42_I8_n331, B1 => mult_42_I8_n332, B2 => 
                           mult_42_I8_n333, ZN => mult_42_I8_n35);
   mult_42_I8_U267 : XOR2_X1 port map( A => B(78), B => x_vector_73_port, Z => 
                           mult_42_I8_n323);
   mult_42_I8_U266 : AOI22_X1 port map( A1 => mult_42_I8_n323, A2 => 
                           mult_42_I8_n318, B1 => mult_42_I8_n319, B2 => 
                           mult_42_I8_n329, ZN => mult_42_I8_n50);
   mult_42_I8_U265 : OAI22_X1 port map( A1 => mult_42_I8_n325, A2 => 
                           mult_42_I8_n326, B1 => mult_42_I8_n327, B2 => 
                           mult_42_I8_n328, ZN => mult_42_I8_n321);
   mult_42_I8_U264 : AOI22_X1 port map( A1 => mult_42_I8_n306, A2 => 
                           mult_42_I8_n318, B1 => mult_42_I8_n319, B2 => 
                           mult_42_I8_n323, ZN => mult_42_I8_n322);
   mult_42_I8_U263 : NAND2_X1 port map( A1 => mult_42_I8_n310, A2 => 
                           mult_42_I8_n322, ZN => mult_42_I8_n57);
   mult_42_I8_U262 : XOR2_X1 port map( A => mult_42_I8_n321, B => 
                           mult_42_I8_n322, Z => mult_42_I8_n58);
   mult_42_I8_U261 : XNOR2_X2 port map( A => x_vector_78_port, B => 
                           x_vector_77_port, ZN => mult_42_I8_n338);
   mult_42_I8_U260 : XNOR2_X2 port map( A => x_vector_76_port, B => 
                           x_vector_75_port, ZN => mult_42_I8_n327);
   mult_42_I8_U259 : XNOR2_X2 port map( A => x_vector_74_port, B => 
                           x_vector_73_port, ZN => mult_42_I8_n332);
   mult_42_I8_U258 : INV_X1 port map( A => B(71), ZN => mult_42_I8_n312);
   mult_42_I8_U257 : INV_X1 port map( A => B(70), ZN => mult_42_I8_n313);
   mult_42_I8_U256 : INV_X1 port map( A => x_vector_73_port, ZN => 
                           mult_42_I8_n317);
   mult_42_I8_U255 : INV_X1 port map( A => x_vector_70_port, ZN => 
                           mult_42_I8_n320);
   mult_42_I8_U254 : INV_X1 port map( A => x_vector_77_port, ZN => 
                           mult_42_I8_n315);
   mult_42_I8_U253 : INV_X1 port map( A => x_vector_75_port, ZN => 
                           mult_42_I8_n316);
   mult_42_I8_U252 : INV_X1 port map( A => x_vector_79_port, ZN => 
                           mult_42_I8_n314);
   mult_42_I8_U251 : INV_X1 port map( A => mult_42_I8_n367, ZN => 
                           mult_42_I8_n298);
   mult_42_I8_U250 : INV_X1 port map( A => mult_42_I8_n374, ZN => 
                           mult_42_I8_n300);
   mult_42_I8_U249 : INV_X1 port map( A => mult_42_I8_n25, ZN => 
                           mult_42_I8_n301);
   mult_42_I8_U248 : INV_X1 port map( A => mult_42_I8_n35, ZN => 
                           mult_42_I8_n299);
   mult_42_I8_U247 : INV_X1 port map( A => mult_42_I8_n90, ZN => 
                           mult_42_I8_n311);
   mult_42_I8_U246 : INV_X1 port map( A => mult_42_I8_n50, ZN => 
                           mult_42_I8_n297);
   mult_42_I8_U245 : INV_X1 port map( A => mult_42_I8_n349, ZN => 
                           mult_42_I8_n295);
   mult_42_I8_U244 : INV_X1 port map( A => mult_42_I8_n383, ZN => 
                           mult_42_I8_n302);
   mult_42_I8_U243 : INV_X1 port map( A => mult_42_I8_n351, ZN => 
                           mult_42_I8_n318);
   mult_42_I8_U242 : INV_X1 port map( A => mult_42_I8_n352, ZN => 
                           mult_42_I8_n319);
   mult_42_I8_U241 : INV_X1 port map( A => mult_42_I8_n324, ZN => 
                           mult_42_I8_n306);
   mult_42_I8_U240 : INV_X1 port map( A => mult_42_I8_n84, ZN => 
                           mult_42_I8_n308);
   mult_42_I8_U239 : INV_X1 port map( A => mult_42_I8_n87, ZN => 
                           mult_42_I8_n309);
   mult_42_I8_U238 : INV_X1 port map( A => mult_42_I8_n321, ZN => 
                           mult_42_I8_n310);
   mult_42_I8_U237 : INV_X1 port map( A => mult_42_I8_n1, ZN => N142);
   mult_42_I8_U236 : INV_X1 port map( A => mult_42_I8_n19, ZN => 
                           mult_42_I8_n303);
   mult_42_I8_U235 : INV_X1 port map( A => mult_42_I8_n74, ZN => 
                           mult_42_I8_n305);
   mult_42_I8_U234 : INV_X1 port map( A => mult_42_I8_n79, ZN => 
                           mult_42_I8_n307);
   mult_42_I8_U233 : INV_X1 port map( A => mult_42_I8_n60, ZN => 
                           mult_42_I8_n296);
   mult_42_I8_U232 : INV_X1 port map( A => mult_42_I8_n67, ZN => 
                           mult_42_I8_n304);
   mult_42_I8_U56 : HA_X1 port map( A => mult_42_I8_n148, B => mult_42_I8_n157,
                           CO => mult_42_I8_n89, S => mult_42_I8_n90);
   mult_42_I8_U55 : FA_X1 port map( A => mult_42_I8_n156, B => mult_42_I8_n139,
                           CI => mult_42_I8_n147, CO => mult_42_I8_n87, S => 
                           mult_42_I8_n88);
   mult_42_I8_U54 : HA_X1 port map( A => mult_42_I8_n107, B => mult_42_I8_n138,
                           CO => mult_42_I8_n85, S => mult_42_I8_n86);
   mult_42_I8_U53 : FA_X1 port map( A => mult_42_I8_n146, B => mult_42_I8_n155,
                           CI => mult_42_I8_n86, CO => mult_42_I8_n83, S => 
                           mult_42_I8_n84);
   mult_42_I8_U52 : FA_X1 port map( A => mult_42_I8_n154, B => mult_42_I8_n129,
                           CI => mult_42_I8_n145, CO => mult_42_I8_n81, S => 
                           mult_42_I8_n82);
   mult_42_I8_U51 : FA_X1 port map( A => mult_42_I8_n85, B => mult_42_I8_n137, 
                           CI => mult_42_I8_n82, CO => mult_42_I8_n79, S => 
                           mult_42_I8_n80);
   mult_42_I8_U50 : HA_X1 port map( A => mult_42_I8_n106, B => mult_42_I8_n128,
                           CO => mult_42_I8_n77, S => mult_42_I8_n78);
   mult_42_I8_U49 : FA_X1 port map( A => mult_42_I8_n136, B => mult_42_I8_n153,
                           CI => mult_42_I8_n144, CO => mult_42_I8_n75, S => 
                           mult_42_I8_n76);
   mult_42_I8_U48 : FA_X1 port map( A => mult_42_I8_n81, B => mult_42_I8_n78, 
                           CI => mult_42_I8_n76, CO => mult_42_I8_n73, S => 
                           mult_42_I8_n74);
   mult_42_I8_U47 : FA_X1 port map( A => mult_42_I8_n135, B => mult_42_I8_n119,
                           CI => mult_42_I8_n152, CO => mult_42_I8_n71, S => 
                           mult_42_I8_n72);
   mult_42_I8_U46 : FA_X1 port map( A => mult_42_I8_n127, B => mult_42_I8_n143,
                           CI => mult_42_I8_n77, CO => mult_42_I8_n69, S => 
                           mult_42_I8_n70);
   mult_42_I8_U45 : FA_X1 port map( A => mult_42_I8_n72, B => mult_42_I8_n75, 
                           CI => mult_42_I8_n70, CO => mult_42_I8_n67, S => 
                           mult_42_I8_n68);
   mult_42_I8_U44 : HA_X1 port map( A => mult_42_I8_n105, B => mult_42_I8_n118,
                           CO => mult_42_I8_n65, S => mult_42_I8_n66);
   mult_42_I8_U43 : FA_X1 port map( A => mult_42_I8_n126, B => mult_42_I8_n134,
                           CI => mult_42_I8_n142, CO => mult_42_I8_n63, S => 
                           mult_42_I8_n64);
   mult_42_I8_U42 : FA_X1 port map( A => mult_42_I8_n66, B => mult_42_I8_n151, 
                           CI => mult_42_I8_n71, CO => mult_42_I8_n61, S => 
                           mult_42_I8_n62);
   mult_42_I8_U41 : FA_X1 port map( A => mult_42_I8_n64, B => mult_42_I8_n69, 
                           CI => mult_42_I8_n62, CO => mult_42_I8_n59, S => 
                           mult_42_I8_n60);
   mult_42_I8_U38 : FA_X1 port map( A => mult_42_I8_n133, B => mult_42_I8_n117,
                           CI => mult_42_I8_n295, CO => mult_42_I8_n55, S => 
                           mult_42_I8_n56);
   mult_42_I8_U37 : FA_X1 port map( A => mult_42_I8_n58, B => mult_42_I8_n65, 
                           CI => mult_42_I8_n63, CO => mult_42_I8_n53, S => 
                           mult_42_I8_n54);
   mult_42_I8_U36 : FA_X1 port map( A => mult_42_I8_n61, B => mult_42_I8_n56, 
                           CI => mult_42_I8_n54, CO => mult_42_I8_n51, S => 
                           mult_42_I8_n52);
   mult_42_I8_U34 : FA_X1 port map( A => mult_42_I8_n124, B => mult_42_I8_n116,
                           CI => mult_42_I8_n132, CO => mult_42_I8_n47, S => 
                           mult_42_I8_n48);
   mult_42_I8_U33 : FA_X1 port map( A => mult_42_I8_n57, B => mult_42_I8_n50, 
                           CI => mult_42_I8_n55, CO => mult_42_I8_n45, S => 
                           mult_42_I8_n46);
   mult_42_I8_U32 : FA_X1 port map( A => mult_42_I8_n53, B => mult_42_I8_n48, 
                           CI => mult_42_I8_n46, CO => mult_42_I8_n43, S => 
                           mult_42_I8_n44);
   mult_42_I8_U31 : FA_X1 port map( A => mult_42_I8_n123, B => mult_42_I8_n115,
                           CI => mult_42_I8_n140, CO => mult_42_I8_n41, S => 
                           mult_42_I8_n42);
   mult_42_I8_U30 : FA_X1 port map( A => mult_42_I8_n297, B => mult_42_I8_n131,
                           CI => mult_42_I8_n47, CO => mult_42_I8_n39, S => 
                           mult_42_I8_n40);
   mult_42_I8_U29 : FA_X1 port map( A => mult_42_I8_n45, B => mult_42_I8_n42, 
                           CI => mult_42_I8_n40, CO => mult_42_I8_n37, S => 
                           mult_42_I8_n38);
   mult_42_I8_U27 : FA_X1 port map( A => mult_42_I8_n114, B => mult_42_I8_n122,
                           CI => mult_42_I8_n299, CO => mult_42_I8_n33, S => 
                           mult_42_I8_n34);
   mult_42_I8_U26 : FA_X1 port map( A => mult_42_I8_n34, B => mult_42_I8_n41, 
                           CI => mult_42_I8_n39, CO => mult_42_I8_n31, S => 
                           mult_42_I8_n32);
   mult_42_I8_U25 : FA_X1 port map( A => mult_42_I8_n121, B => mult_42_I8_n35, 
                           CI => mult_42_I8_n298, CO => mult_42_I8_n29, S => 
                           mult_42_I8_n30);
   mult_42_I8_U24 : FA_X1 port map( A => mult_42_I8_n33, B => mult_42_I8_n113, 
                           CI => mult_42_I8_n30, CO => mult_42_I8_n27, S => 
                           mult_42_I8_n28);
   mult_42_I8_U22 : FA_X1 port map( A => mult_42_I8_n301, B => mult_42_I8_n112,
                           CI => mult_42_I8_n29, CO => mult_42_I8_n23, S => 
                           mult_42_I8_n24);
   mult_42_I8_U21 : FA_X1 port map( A => mult_42_I8_n111, B => mult_42_I8_n25, 
                           CI => mult_42_I8_n300, CO => mult_42_I8_n21, S => 
                           mult_42_I8_n22);
   mult_42_I8_U10 : FA_X1 port map( A => mult_42_I8_n52, B => mult_42_I8_n59, 
                           CI => mult_42_I8_n10, CO => mult_42_I8_n9, S => N133
                           );
   mult_42_I8_U9 : FA_X1 port map( A => mult_42_I8_n44, B => mult_42_I8_n51, CI
                           => mult_42_I8_n9, CO => mult_42_I8_n8, S => N134);
   mult_42_I8_U8 : FA_X1 port map( A => mult_42_I8_n38, B => mult_42_I8_n43, CI
                           => mult_42_I8_n8, CO => mult_42_I8_n7, S => N135);
   mult_42_I8_U7 : FA_X1 port map( A => mult_42_I8_n32, B => mult_42_I8_n37, CI
                           => mult_42_I8_n7, CO => mult_42_I8_n6, S => N136);
   mult_42_I8_U6 : FA_X1 port map( A => mult_42_I8_n28, B => mult_42_I8_n31, CI
                           => mult_42_I8_n6, CO => mult_42_I8_n5, S => N137);
   mult_42_I8_U5 : FA_X1 port map( A => mult_42_I8_n24, B => mult_42_I8_n27, CI
                           => mult_42_I8_n5, CO => mult_42_I8_n4, S => N138);
   mult_42_I8_U4 : FA_X1 port map( A => mult_42_I8_n23, B => mult_42_I8_n22, CI
                           => mult_42_I8_n4, CO => mult_42_I8_n3, S => N139);
   mult_42_I8_U3 : FA_X1 port map( A => mult_42_I8_n21, B => mult_42_I8_n303, 
                           CI => mult_42_I8_n3, CO => mult_42_I8_n2, S => N140)
                           ;
   mult_42_I8_U2 : FA_X1 port map( A => mult_42_I8_n302, B => mult_42_I8_n19, 
                           CI => mult_42_I8_n2, CO => mult_42_I8_n1, S => N141)
                           ;
   mult_42_I9_U391 : NAND2_X1 port map( A1 => x_vector_81_port, A2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n341);
   mult_42_I9_U390 : XNOR2_X1 port map( A => B(82), B => x_vector_81_port, ZN 
                           => mult_42_I9_n340);
   mult_42_I9_U389 : OAI22_X1 port map( A1 => B(81), A2 => mult_42_I9_n341, B1 
                           => mult_42_I9_n340, B2 => mult_42_I9_n320, ZN => 
                           mult_42_I9_n402);
   mult_42_I9_U388 : NAND3_X1 port map( A1 => mult_42_I9_n402, A2 => 
                           mult_42_I9_n312, A3 => x_vector_81_port, ZN => 
                           mult_42_I9_n400);
   mult_42_I9_U387 : XNOR2_X1 port map( A => x_vector_82_port, B => 
                           x_vector_81_port, ZN => mult_42_I9_n352);
   mult_42_I9_U386 : NAND2_X1 port map( A1 => mult_42_I9_n319, A2 => 
                           mult_42_I9_n402, ZN => mult_42_I9_n401);
   mult_42_I9_U385 : MUX2_X1 port map( A => mult_42_I9_n400, B => 
                           mult_42_I9_n401, S => B(80), Z => mult_42_I9_n396);
   mult_42_I9_U384 : XOR2_X1 port map( A => x_vector_83_port, B => 
                           x_vector_82_port, Z => mult_42_I9_n399);
   mult_42_I9_U383 : NAND2_X1 port map( A1 => mult_42_I9_n352, A2 => 
                           mult_42_I9_n399, ZN => mult_42_I9_n351);
   mult_42_I9_U382 : NOR3_X1 port map( A1 => mult_42_I9_n352, A2 => B(80), A3 
                           => mult_42_I9_n317, ZN => mult_42_I9_n398);
   mult_42_I9_U381 : AOI21_X1 port map( B1 => x_vector_83_port, B2 => 
                           mult_42_I9_n318, A => mult_42_I9_n398, ZN => 
                           mult_42_I9_n397);
   mult_42_I9_U380 : OAI222_X1 port map( A1 => mult_42_I9_n396, A2 => 
                           mult_42_I9_n311, B1 => mult_42_I9_n397, B2 => 
                           mult_42_I9_n396, C1 => mult_42_I9_n397, C2 => 
                           mult_42_I9_n311, ZN => mult_42_I9_n395);
   mult_42_I9_U379 : AOI222_X1 port map( A1 => mult_42_I9_n395, A2 => 
                           mult_42_I9_n88, B1 => mult_42_I9_n395, B2 => 
                           mult_42_I9_n89, C1 => mult_42_I9_n89, C2 => 
                           mult_42_I9_n88, ZN => mult_42_I9_n394);
   mult_42_I9_U378 : OAI222_X1 port map( A1 => mult_42_I9_n394, A2 => 
                           mult_42_I9_n308, B1 => mult_42_I9_n394, B2 => 
                           mult_42_I9_n309, C1 => mult_42_I9_n309, C2 => 
                           mult_42_I9_n308, ZN => mult_42_I9_n393);
   mult_42_I9_U377 : AOI222_X1 port map( A1 => mult_42_I9_n393, A2 => 
                           mult_42_I9_n80, B1 => mult_42_I9_n393, B2 => 
                           mult_42_I9_n83, C1 => mult_42_I9_n83, C2 => 
                           mult_42_I9_n80, ZN => mult_42_I9_n392);
   mult_42_I9_U376 : OAI222_X1 port map( A1 => mult_42_I9_n392, A2 => 
                           mult_42_I9_n305, B1 => mult_42_I9_n392, B2 => 
                           mult_42_I9_n307, C1 => mult_42_I9_n307, C2 => 
                           mult_42_I9_n305, ZN => mult_42_I9_n391);
   mult_42_I9_U375 : AOI222_X1 port map( A1 => mult_42_I9_n391, A2 => 
                           mult_42_I9_n68, B1 => mult_42_I9_n391, B2 => 
                           mult_42_I9_n73, C1 => mult_42_I9_n73, C2 => 
                           mult_42_I9_n68, ZN => mult_42_I9_n390);
   mult_42_I9_U374 : OAI222_X1 port map( A1 => mult_42_I9_n390, A2 => 
                           mult_42_I9_n296, B1 => mult_42_I9_n390, B2 => 
                           mult_42_I9_n304, C1 => mult_42_I9_n304, C2 => 
                           mult_42_I9_n296, ZN => mult_42_I9_n10);
   mult_42_I9_U373 : XOR2_X1 port map( A => x_vector_89_port, B => 
                           x_vector_88_port, Z => mult_42_I9_n389);
   mult_42_I9_U372 : NAND2_X1 port map( A1 => mult_42_I9_n338, A2 => 
                           mult_42_I9_n389, ZN => mult_42_I9_n337);
   mult_42_I9_U371 : OR3_X1 port map( A1 => mult_42_I9_n338, A2 => B(80), A3 =>
                           mult_42_I9_n314, ZN => mult_42_I9_n388);
   mult_42_I9_U370 : OAI21_X1 port map( B1 => mult_42_I9_n314, B2 => 
                           mult_42_I9_n337, A => mult_42_I9_n388, ZN => 
                           mult_42_I9_n105);
   mult_42_I9_U369 : XOR2_X1 port map( A => x_vector_87_port, B => 
                           x_vector_86_port, Z => mult_42_I9_n387);
   mult_42_I9_U368 : NAND2_X1 port map( A1 => mult_42_I9_n327, A2 => 
                           mult_42_I9_n387, ZN => mult_42_I9_n326);
   mult_42_I9_U367 : OR3_X1 port map( A1 => mult_42_I9_n327, A2 => B(80), A3 =>
                           mult_42_I9_n315, ZN => mult_42_I9_n386);
   mult_42_I9_U366 : OAI21_X1 port map( B1 => mult_42_I9_n315, B2 => 
                           mult_42_I9_n326, A => mult_42_I9_n386, ZN => 
                           mult_42_I9_n106);
   mult_42_I9_U365 : XOR2_X1 port map( A => x_vector_85_port, B => 
                           x_vector_84_port, Z => mult_42_I9_n385);
   mult_42_I9_U364 : NAND2_X1 port map( A1 => mult_42_I9_n332, A2 => 
                           mult_42_I9_n385, ZN => mult_42_I9_n331);
   mult_42_I9_U363 : OR3_X1 port map( A1 => mult_42_I9_n332, A2 => B(80), A3 =>
                           mult_42_I9_n316, ZN => mult_42_I9_n384);
   mult_42_I9_U362 : OAI21_X1 port map( B1 => mult_42_I9_n316, B2 => 
                           mult_42_I9_n331, A => mult_42_I9_n384, ZN => 
                           mult_42_I9_n107);
   mult_42_I9_U361 : XOR2_X1 port map( A => B(89), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n339);
   mult_42_I9_U360 : OAI22_X1 port map( A1 => mult_42_I9_n339, A2 => 
                           mult_42_I9_n338, B1 => mult_42_I9_n337, B2 => 
                           mult_42_I9_n339, ZN => mult_42_I9_n383);
   mult_42_I9_U359 : XOR2_X1 port map( A => B(87), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n382);
   mult_42_I9_U358 : XOR2_X1 port map( A => B(88), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n336);
   mult_42_I9_U357 : OAI22_X1 port map( A1 => mult_42_I9_n382, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n336, ZN => mult_42_I9_n111);
   mult_42_I9_U356 : XOR2_X1 port map( A => B(86), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n381);
   mult_42_I9_U355 : OAI22_X1 port map( A1 => mult_42_I9_n381, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n382, ZN => mult_42_I9_n112);
   mult_42_I9_U354 : XOR2_X1 port map( A => B(85), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n380);
   mult_42_I9_U353 : OAI22_X1 port map( A1 => mult_42_I9_n380, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n381, ZN => mult_42_I9_n113);
   mult_42_I9_U352 : XOR2_X1 port map( A => B(84), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n379);
   mult_42_I9_U351 : OAI22_X1 port map( A1 => mult_42_I9_n379, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n380, ZN => mult_42_I9_n114);
   mult_42_I9_U350 : XOR2_X1 port map( A => B(83), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n378);
   mult_42_I9_U349 : OAI22_X1 port map( A1 => mult_42_I9_n378, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n379, ZN => mult_42_I9_n115);
   mult_42_I9_U348 : XOR2_X1 port map( A => B(82), B => mult_42_I9_n314, Z => 
                           mult_42_I9_n377);
   mult_42_I9_U347 : OAI22_X1 port map( A1 => mult_42_I9_n377, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n378, ZN => mult_42_I9_n116);
   mult_42_I9_U346 : XOR2_X1 port map( A => mult_42_I9_n312, B => 
                           x_vector_89_port, Z => mult_42_I9_n376);
   mult_42_I9_U345 : OAI22_X1 port map( A1 => mult_42_I9_n376, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n377, ZN => mult_42_I9_n117);
   mult_42_I9_U344 : XOR2_X1 port map( A => mult_42_I9_n314, B => B(80), Z => 
                           mult_42_I9_n375);
   mult_42_I9_U343 : OAI22_X1 port map( A1 => mult_42_I9_n375, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n376, ZN => mult_42_I9_n118);
   mult_42_I9_U342 : NOR2_X1 port map( A1 => mult_42_I9_n338, A2 => 
                           mult_42_I9_n313, ZN => mult_42_I9_n119);
   mult_42_I9_U341 : XOR2_X1 port map( A => B(89), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n335);
   mult_42_I9_U340 : OAI22_X1 port map( A1 => mult_42_I9_n335, A2 => 
                           mult_42_I9_n327, B1 => mult_42_I9_n326, B2 => 
                           mult_42_I9_n335, ZN => mult_42_I9_n374);
   mult_42_I9_U339 : XOR2_X1 port map( A => B(87), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n373);
   mult_42_I9_U338 : XOR2_X1 port map( A => B(88), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n334);
   mult_42_I9_U337 : OAI22_X1 port map( A1 => mult_42_I9_n373, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n334, ZN => mult_42_I9_n121);
   mult_42_I9_U336 : XOR2_X1 port map( A => B(86), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n372);
   mult_42_I9_U335 : OAI22_X1 port map( A1 => mult_42_I9_n372, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n373, ZN => mult_42_I9_n122);
   mult_42_I9_U334 : XOR2_X1 port map( A => B(85), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n371);
   mult_42_I9_U333 : OAI22_X1 port map( A1 => mult_42_I9_n371, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n372, ZN => mult_42_I9_n123);
   mult_42_I9_U332 : XOR2_X1 port map( A => B(84), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n328);
   mult_42_I9_U331 : OAI22_X1 port map( A1 => mult_42_I9_n328, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n371, ZN => mult_42_I9_n124);
   mult_42_I9_U330 : XOR2_X1 port map( A => B(82), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n370);
   mult_42_I9_U329 : XOR2_X1 port map( A => B(83), B => mult_42_I9_n315, Z => 
                           mult_42_I9_n325);
   mult_42_I9_U328 : OAI22_X1 port map( A1 => mult_42_I9_n370, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n325, ZN => mult_42_I9_n126);
   mult_42_I9_U327 : XOR2_X1 port map( A => mult_42_I9_n312, B => 
                           x_vector_87_port, Z => mult_42_I9_n369);
   mult_42_I9_U326 : OAI22_X1 port map( A1 => mult_42_I9_n369, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n370, ZN => mult_42_I9_n127);
   mult_42_I9_U325 : XOR2_X1 port map( A => mult_42_I9_n313, B => 
                           x_vector_87_port, Z => mult_42_I9_n368);
   mult_42_I9_U324 : OAI22_X1 port map( A1 => mult_42_I9_n368, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n369, ZN => mult_42_I9_n128);
   mult_42_I9_U323 : NOR2_X1 port map( A1 => mult_42_I9_n327, A2 => 
                           mult_42_I9_n313, ZN => mult_42_I9_n129);
   mult_42_I9_U322 : XOR2_X1 port map( A => B(89), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n333);
   mult_42_I9_U321 : OAI22_X1 port map( A1 => mult_42_I9_n333, A2 => 
                           mult_42_I9_n332, B1 => mult_42_I9_n331, B2 => 
                           mult_42_I9_n333, ZN => mult_42_I9_n367);
   mult_42_I9_U320 : XOR2_X1 port map( A => B(87), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n366);
   mult_42_I9_U319 : XOR2_X1 port map( A => B(88), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n330);
   mult_42_I9_U318 : OAI22_X1 port map( A1 => mult_42_I9_n366, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n330, ZN => mult_42_I9_n131);
   mult_42_I9_U317 : XOR2_X1 port map( A => B(86), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n365);
   mult_42_I9_U316 : OAI22_X1 port map( A1 => mult_42_I9_n365, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n366, ZN => mult_42_I9_n132);
   mult_42_I9_U315 : XOR2_X1 port map( A => B(85), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n364);
   mult_42_I9_U314 : OAI22_X1 port map( A1 => mult_42_I9_n364, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n365, ZN => mult_42_I9_n133);
   mult_42_I9_U313 : XOR2_X1 port map( A => B(84), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n363);
   mult_42_I9_U312 : OAI22_X1 port map( A1 => mult_42_I9_n363, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n364, ZN => mult_42_I9_n134);
   mult_42_I9_U311 : XOR2_X1 port map( A => B(83), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n362);
   mult_42_I9_U310 : OAI22_X1 port map( A1 => mult_42_I9_n362, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n363, ZN => mult_42_I9_n135);
   mult_42_I9_U309 : XOR2_X1 port map( A => B(82), B => mult_42_I9_n316, Z => 
                           mult_42_I9_n361);
   mult_42_I9_U308 : OAI22_X1 port map( A1 => mult_42_I9_n361, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n362, ZN => mult_42_I9_n136);
   mult_42_I9_U307 : XOR2_X1 port map( A => mult_42_I9_n312, B => 
                           x_vector_85_port, Z => mult_42_I9_n360);
   mult_42_I9_U306 : OAI22_X1 port map( A1 => mult_42_I9_n360, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n361, ZN => mult_42_I9_n137);
   mult_42_I9_U305 : XOR2_X1 port map( A => mult_42_I9_n313, B => 
                           x_vector_85_port, Z => mult_42_I9_n359);
   mult_42_I9_U304 : OAI22_X1 port map( A1 => mult_42_I9_n359, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n360, ZN => mult_42_I9_n138);
   mult_42_I9_U303 : NOR2_X1 port map( A1 => mult_42_I9_n332, A2 => 
                           mult_42_I9_n313, ZN => mult_42_I9_n139);
   mult_42_I9_U302 : XOR2_X1 port map( A => B(89), B => x_vector_83_port, Z => 
                           mult_42_I9_n329);
   mult_42_I9_U301 : AOI22_X1 port map( A1 => mult_42_I9_n329, A2 => 
                           mult_42_I9_n319, B1 => mult_42_I9_n318, B2 => 
                           mult_42_I9_n329, ZN => mult_42_I9_n140);
   mult_42_I9_U300 : XOR2_X1 port map( A => B(86), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n358);
   mult_42_I9_U299 : XOR2_X1 port map( A => B(87), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n324);
   mult_42_I9_U298 : OAI22_X1 port map( A1 => mult_42_I9_n358, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n324, ZN => mult_42_I9_n142);
   mult_42_I9_U297 : XOR2_X1 port map( A => B(85), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n357);
   mult_42_I9_U296 : OAI22_X1 port map( A1 => mult_42_I9_n357, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n358, ZN => mult_42_I9_n143);
   mult_42_I9_U295 : XOR2_X1 port map( A => B(84), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n356);
   mult_42_I9_U294 : OAI22_X1 port map( A1 => mult_42_I9_n356, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n357, ZN => mult_42_I9_n144);
   mult_42_I9_U293 : XOR2_X1 port map( A => B(83), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n355);
   mult_42_I9_U292 : OAI22_X1 port map( A1 => mult_42_I9_n355, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n356, ZN => mult_42_I9_n145);
   mult_42_I9_U291 : XOR2_X1 port map( A => B(82), B => mult_42_I9_n317, Z => 
                           mult_42_I9_n354);
   mult_42_I9_U290 : OAI22_X1 port map( A1 => mult_42_I9_n354, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n355, ZN => mult_42_I9_n146);
   mult_42_I9_U289 : XOR2_X1 port map( A => mult_42_I9_n312, B => 
                           x_vector_83_port, Z => mult_42_I9_n353);
   mult_42_I9_U288 : OAI22_X1 port map( A1 => mult_42_I9_n353, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n354, ZN => mult_42_I9_n147);
   mult_42_I9_U287 : XOR2_X1 port map( A => mult_42_I9_n313, B => 
                           x_vector_83_port, Z => mult_42_I9_n350);
   mult_42_I9_U286 : OAI22_X1 port map( A1 => mult_42_I9_n350, A2 => 
                           mult_42_I9_n351, B1 => mult_42_I9_n352, B2 => 
                           mult_42_I9_n353, ZN => mult_42_I9_n148);
   mult_42_I9_U285 : XNOR2_X1 port map( A => B(89), B => x_vector_81_port, ZN 
                           => mult_42_I9_n348);
   mult_42_I9_U284 : OAI22_X1 port map( A1 => mult_42_I9_n320, A2 => 
                           mult_42_I9_n348, B1 => mult_42_I9_n341, B2 => 
                           mult_42_I9_n348, ZN => mult_42_I9_n349);
   mult_42_I9_U283 : XNOR2_X1 port map( A => B(88), B => x_vector_81_port, ZN 
                           => mult_42_I9_n347);
   mult_42_I9_U282 : OAI22_X1 port map( A1 => mult_42_I9_n347, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n348, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n151);
   mult_42_I9_U281 : XNOR2_X1 port map( A => B(87), B => x_vector_81_port, ZN 
                           => mult_42_I9_n346);
   mult_42_I9_U280 : OAI22_X1 port map( A1 => mult_42_I9_n346, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n347, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n152);
   mult_42_I9_U279 : XNOR2_X1 port map( A => B(86), B => x_vector_81_port, ZN 
                           => mult_42_I9_n345);
   mult_42_I9_U278 : OAI22_X1 port map( A1 => mult_42_I9_n345, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n346, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n153);
   mult_42_I9_U277 : XNOR2_X1 port map( A => B(85), B => x_vector_81_port, ZN 
                           => mult_42_I9_n344);
   mult_42_I9_U276 : OAI22_X1 port map( A1 => mult_42_I9_n344, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n345, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n154);
   mult_42_I9_U275 : XNOR2_X1 port map( A => B(84), B => x_vector_81_port, ZN 
                           => mult_42_I9_n343);
   mult_42_I9_U274 : OAI22_X1 port map( A1 => mult_42_I9_n343, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n344, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n155);
   mult_42_I9_U273 : XNOR2_X1 port map( A => B(83), B => x_vector_81_port, ZN 
                           => mult_42_I9_n342);
   mult_42_I9_U272 : OAI22_X1 port map( A1 => mult_42_I9_n342, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n343, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n156);
   mult_42_I9_U271 : OAI22_X1 port map( A1 => mult_42_I9_n340, A2 => 
                           mult_42_I9_n341, B1 => mult_42_I9_n342, B2 => 
                           mult_42_I9_n320, ZN => mult_42_I9_n157);
   mult_42_I9_U270 : OAI22_X1 port map( A1 => mult_42_I9_n336, A2 => 
                           mult_42_I9_n337, B1 => mult_42_I9_n338, B2 => 
                           mult_42_I9_n339, ZN => mult_42_I9_n19);
   mult_42_I9_U269 : OAI22_X1 port map( A1 => mult_42_I9_n334, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n335, ZN => mult_42_I9_n25);
   mult_42_I9_U268 : OAI22_X1 port map( A1 => mult_42_I9_n330, A2 => 
                           mult_42_I9_n331, B1 => mult_42_I9_n332, B2 => 
                           mult_42_I9_n333, ZN => mult_42_I9_n35);
   mult_42_I9_U267 : XOR2_X1 port map( A => B(88), B => x_vector_83_port, Z => 
                           mult_42_I9_n323);
   mult_42_I9_U266 : AOI22_X1 port map( A1 => mult_42_I9_n323, A2 => 
                           mult_42_I9_n318, B1 => mult_42_I9_n319, B2 => 
                           mult_42_I9_n329, ZN => mult_42_I9_n50);
   mult_42_I9_U265 : OAI22_X1 port map( A1 => mult_42_I9_n325, A2 => 
                           mult_42_I9_n326, B1 => mult_42_I9_n327, B2 => 
                           mult_42_I9_n328, ZN => mult_42_I9_n321);
   mult_42_I9_U264 : AOI22_X1 port map( A1 => mult_42_I9_n306, A2 => 
                           mult_42_I9_n318, B1 => mult_42_I9_n319, B2 => 
                           mult_42_I9_n323, ZN => mult_42_I9_n322);
   mult_42_I9_U263 : NAND2_X1 port map( A1 => mult_42_I9_n310, A2 => 
                           mult_42_I9_n322, ZN => mult_42_I9_n57);
   mult_42_I9_U262 : XOR2_X1 port map( A => mult_42_I9_n321, B => 
                           mult_42_I9_n322, Z => mult_42_I9_n58);
   mult_42_I9_U261 : XNOR2_X2 port map( A => x_vector_88_port, B => 
                           x_vector_87_port, ZN => mult_42_I9_n338);
   mult_42_I9_U260 : XNOR2_X2 port map( A => x_vector_86_port, B => 
                           x_vector_85_port, ZN => mult_42_I9_n327);
   mult_42_I9_U259 : XNOR2_X2 port map( A => x_vector_84_port, B => 
                           x_vector_83_port, ZN => mult_42_I9_n332);
   mult_42_I9_U258 : INV_X1 port map( A => B(81), ZN => mult_42_I9_n312);
   mult_42_I9_U257 : INV_X1 port map( A => B(80), ZN => mult_42_I9_n313);
   mult_42_I9_U256 : INV_X1 port map( A => x_vector_83_port, ZN => 
                           mult_42_I9_n317);
   mult_42_I9_U255 : INV_X1 port map( A => x_vector_80_port, ZN => 
                           mult_42_I9_n320);
   mult_42_I9_U254 : INV_X1 port map( A => x_vector_87_port, ZN => 
                           mult_42_I9_n315);
   mult_42_I9_U253 : INV_X1 port map( A => x_vector_85_port, ZN => 
                           mult_42_I9_n316);
   mult_42_I9_U252 : INV_X1 port map( A => x_vector_89_port, ZN => 
                           mult_42_I9_n314);
   mult_42_I9_U251 : INV_X1 port map( A => mult_42_I9_n374, ZN => 
                           mult_42_I9_n300);
   mult_42_I9_U250 : INV_X1 port map( A => mult_42_I9_n25, ZN => 
                           mult_42_I9_n301);
   mult_42_I9_U249 : INV_X1 port map( A => mult_42_I9_n90, ZN => 
                           mult_42_I9_n311);
   mult_42_I9_U248 : INV_X1 port map( A => mult_42_I9_n50, ZN => 
                           mult_42_I9_n297);
   mult_42_I9_U247 : INV_X1 port map( A => mult_42_I9_n367, ZN => 
                           mult_42_I9_n298);
   mult_42_I9_U246 : INV_X1 port map( A => mult_42_I9_n349, ZN => 
                           mult_42_I9_n295);
   mult_42_I9_U245 : INV_X1 port map( A => mult_42_I9_n383, ZN => 
                           mult_42_I9_n302);
   mult_42_I9_U244 : INV_X1 port map( A => mult_42_I9_n35, ZN => 
                           mult_42_I9_n299);
   mult_42_I9_U243 : INV_X1 port map( A => mult_42_I9_n351, ZN => 
                           mult_42_I9_n318);
   mult_42_I9_U242 : INV_X1 port map( A => mult_42_I9_n352, ZN => 
                           mult_42_I9_n319);
   mult_42_I9_U241 : INV_X1 port map( A => mult_42_I9_n324, ZN => 
                           mult_42_I9_n306);
   mult_42_I9_U240 : INV_X1 port map( A => mult_42_I9_n84, ZN => 
                           mult_42_I9_n308);
   mult_42_I9_U239 : INV_X1 port map( A => mult_42_I9_n87, ZN => 
                           mult_42_I9_n309);
   mult_42_I9_U238 : INV_X1 port map( A => mult_42_I9_n19, ZN => 
                           mult_42_I9_n303);
   mult_42_I9_U237 : INV_X1 port map( A => mult_42_I9_n321, ZN => 
                           mult_42_I9_n310);
   mult_42_I9_U236 : INV_X1 port map( A => mult_42_I9_n1, ZN => N162_port);
   mult_42_I9_U235 : INV_X1 port map( A => mult_42_I9_n74, ZN => 
                           mult_42_I9_n305);
   mult_42_I9_U234 : INV_X1 port map( A => mult_42_I9_n79, ZN => 
                           mult_42_I9_n307);
   mult_42_I9_U233 : INV_X1 port map( A => mult_42_I9_n60, ZN => 
                           mult_42_I9_n296);
   mult_42_I9_U232 : INV_X1 port map( A => mult_42_I9_n67, ZN => 
                           mult_42_I9_n304);
   mult_42_I9_U56 : HA_X1 port map( A => mult_42_I9_n148, B => mult_42_I9_n157,
                           CO => mult_42_I9_n89, S => mult_42_I9_n90);
   mult_42_I9_U55 : FA_X1 port map( A => mult_42_I9_n156, B => mult_42_I9_n139,
                           CI => mult_42_I9_n147, CO => mult_42_I9_n87, S => 
                           mult_42_I9_n88);
   mult_42_I9_U54 : HA_X1 port map( A => mult_42_I9_n107, B => mult_42_I9_n138,
                           CO => mult_42_I9_n85, S => mult_42_I9_n86);
   mult_42_I9_U53 : FA_X1 port map( A => mult_42_I9_n146, B => mult_42_I9_n155,
                           CI => mult_42_I9_n86, CO => mult_42_I9_n83, S => 
                           mult_42_I9_n84);
   mult_42_I9_U52 : FA_X1 port map( A => mult_42_I9_n154, B => mult_42_I9_n129,
                           CI => mult_42_I9_n145, CO => mult_42_I9_n81, S => 
                           mult_42_I9_n82);
   mult_42_I9_U51 : FA_X1 port map( A => mult_42_I9_n85, B => mult_42_I9_n137, 
                           CI => mult_42_I9_n82, CO => mult_42_I9_n79, S => 
                           mult_42_I9_n80);
   mult_42_I9_U50 : HA_X1 port map( A => mult_42_I9_n106, B => mult_42_I9_n128,
                           CO => mult_42_I9_n77, S => mult_42_I9_n78);
   mult_42_I9_U49 : FA_X1 port map( A => mult_42_I9_n136, B => mult_42_I9_n153,
                           CI => mult_42_I9_n144, CO => mult_42_I9_n75, S => 
                           mult_42_I9_n76);
   mult_42_I9_U48 : FA_X1 port map( A => mult_42_I9_n81, B => mult_42_I9_n78, 
                           CI => mult_42_I9_n76, CO => mult_42_I9_n73, S => 
                           mult_42_I9_n74);
   mult_42_I9_U47 : FA_X1 port map( A => mult_42_I9_n135, B => mult_42_I9_n119,
                           CI => mult_42_I9_n152, CO => mult_42_I9_n71, S => 
                           mult_42_I9_n72);
   mult_42_I9_U46 : FA_X1 port map( A => mult_42_I9_n127, B => mult_42_I9_n143,
                           CI => mult_42_I9_n77, CO => mult_42_I9_n69, S => 
                           mult_42_I9_n70);
   mult_42_I9_U45 : FA_X1 port map( A => mult_42_I9_n72, B => mult_42_I9_n75, 
                           CI => mult_42_I9_n70, CO => mult_42_I9_n67, S => 
                           mult_42_I9_n68);
   mult_42_I9_U44 : HA_X1 port map( A => mult_42_I9_n105, B => mult_42_I9_n118,
                           CO => mult_42_I9_n65, S => mult_42_I9_n66);
   mult_42_I9_U43 : FA_X1 port map( A => mult_42_I9_n126, B => mult_42_I9_n134,
                           CI => mult_42_I9_n142, CO => mult_42_I9_n63, S => 
                           mult_42_I9_n64);
   mult_42_I9_U42 : FA_X1 port map( A => mult_42_I9_n66, B => mult_42_I9_n151, 
                           CI => mult_42_I9_n71, CO => mult_42_I9_n61, S => 
                           mult_42_I9_n62);
   mult_42_I9_U41 : FA_X1 port map( A => mult_42_I9_n64, B => mult_42_I9_n69, 
                           CI => mult_42_I9_n62, CO => mult_42_I9_n59, S => 
                           mult_42_I9_n60);
   mult_42_I9_U38 : FA_X1 port map( A => mult_42_I9_n133, B => mult_42_I9_n117,
                           CI => mult_42_I9_n295, CO => mult_42_I9_n55, S => 
                           mult_42_I9_n56);
   mult_42_I9_U37 : FA_X1 port map( A => mult_42_I9_n58, B => mult_42_I9_n65, 
                           CI => mult_42_I9_n63, CO => mult_42_I9_n53, S => 
                           mult_42_I9_n54);
   mult_42_I9_U36 : FA_X1 port map( A => mult_42_I9_n61, B => mult_42_I9_n56, 
                           CI => mult_42_I9_n54, CO => mult_42_I9_n51, S => 
                           mult_42_I9_n52);
   mult_42_I9_U34 : FA_X1 port map( A => mult_42_I9_n124, B => mult_42_I9_n116,
                           CI => mult_42_I9_n132, CO => mult_42_I9_n47, S => 
                           mult_42_I9_n48);
   mult_42_I9_U33 : FA_X1 port map( A => mult_42_I9_n57, B => mult_42_I9_n50, 
                           CI => mult_42_I9_n55, CO => mult_42_I9_n45, S => 
                           mult_42_I9_n46);
   mult_42_I9_U32 : FA_X1 port map( A => mult_42_I9_n53, B => mult_42_I9_n48, 
                           CI => mult_42_I9_n46, CO => mult_42_I9_n43, S => 
                           mult_42_I9_n44);
   mult_42_I9_U31 : FA_X1 port map( A => mult_42_I9_n123, B => mult_42_I9_n115,
                           CI => mult_42_I9_n140, CO => mult_42_I9_n41, S => 
                           mult_42_I9_n42);
   mult_42_I9_U30 : FA_X1 port map( A => mult_42_I9_n297, B => mult_42_I9_n131,
                           CI => mult_42_I9_n47, CO => mult_42_I9_n39, S => 
                           mult_42_I9_n40);
   mult_42_I9_U29 : FA_X1 port map( A => mult_42_I9_n45, B => mult_42_I9_n42, 
                           CI => mult_42_I9_n40, CO => mult_42_I9_n37, S => 
                           mult_42_I9_n38);
   mult_42_I9_U27 : FA_X1 port map( A => mult_42_I9_n114, B => mult_42_I9_n122,
                           CI => mult_42_I9_n299, CO => mult_42_I9_n33, S => 
                           mult_42_I9_n34);
   mult_42_I9_U26 : FA_X1 port map( A => mult_42_I9_n34, B => mult_42_I9_n41, 
                           CI => mult_42_I9_n39, CO => mult_42_I9_n31, S => 
                           mult_42_I9_n32);
   mult_42_I9_U25 : FA_X1 port map( A => mult_42_I9_n121, B => mult_42_I9_n35, 
                           CI => mult_42_I9_n298, CO => mult_42_I9_n29, S => 
                           mult_42_I9_n30);
   mult_42_I9_U24 : FA_X1 port map( A => mult_42_I9_n33, B => mult_42_I9_n113, 
                           CI => mult_42_I9_n30, CO => mult_42_I9_n27, S => 
                           mult_42_I9_n28);
   mult_42_I9_U22 : FA_X1 port map( A => mult_42_I9_n301, B => mult_42_I9_n112,
                           CI => mult_42_I9_n29, CO => mult_42_I9_n23, S => 
                           mult_42_I9_n24);
   mult_42_I9_U21 : FA_X1 port map( A => mult_42_I9_n111, B => mult_42_I9_n25, 
                           CI => mult_42_I9_n300, CO => mult_42_I9_n21, S => 
                           mult_42_I9_n22);
   mult_42_I9_U10 : FA_X1 port map( A => mult_42_I9_n52, B => mult_42_I9_n59, 
                           CI => mult_42_I9_n10, CO => mult_42_I9_n9, S => N153
                           );
   mult_42_I9_U9 : FA_X1 port map( A => mult_42_I9_n44, B => mult_42_I9_n51, CI
                           => mult_42_I9_n9, CO => mult_42_I9_n8, S => N154);
   mult_42_I9_U8 : FA_X1 port map( A => mult_42_I9_n38, B => mult_42_I9_n43, CI
                           => mult_42_I9_n8, CO => mult_42_I9_n7, S => N155);
   mult_42_I9_U7 : FA_X1 port map( A => mult_42_I9_n32, B => mult_42_I9_n37, CI
                           => mult_42_I9_n7, CO => mult_42_I9_n6, S => 
                           N156_port);
   mult_42_I9_U6 : FA_X1 port map( A => mult_42_I9_n28, B => mult_42_I9_n31, CI
                           => mult_42_I9_n6, CO => mult_42_I9_n5, S => 
                           N157_port);
   mult_42_I9_U5 : FA_X1 port map( A => mult_42_I9_n24, B => mult_42_I9_n27, CI
                           => mult_42_I9_n5, CO => mult_42_I9_n4, S => 
                           N158_port);
   mult_42_I9_U4 : FA_X1 port map( A => mult_42_I9_n23, B => mult_42_I9_n22, CI
                           => mult_42_I9_n4, CO => mult_42_I9_n3, S => 
                           N159_port);
   mult_42_I9_U3 : FA_X1 port map( A => mult_42_I9_n21, B => mult_42_I9_n303, 
                           CI => mult_42_I9_n3, CO => mult_42_I9_n2, S => 
                           N160_port);
   mult_42_I9_U2 : FA_X1 port map( A => mult_42_I9_n302, B => mult_42_I9_n19, 
                           CI => mult_42_I9_n2, CO => mult_42_I9_n1, S => 
                           N161_port);
   mult_42_I10_U391 : NAND2_X1 port map( A1 => x_vector_91_port, A2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n341);
   mult_42_I10_U390 : XNOR2_X1 port map( A => B(92), B => x_vector_91_port, ZN 
                           => mult_42_I10_n340);
   mult_42_I10_U389 : OAI22_X1 port map( A1 => B(91), A2 => mult_42_I10_n341, 
                           B1 => mult_42_I10_n340, B2 => mult_42_I10_n320, ZN 
                           => mult_42_I10_n402);
   mult_42_I10_U388 : NAND3_X1 port map( A1 => mult_42_I10_n402, A2 => 
                           mult_42_I10_n312, A3 => x_vector_91_port, ZN => 
                           mult_42_I10_n400);
   mult_42_I10_U387 : XNOR2_X1 port map( A => x_vector_92_port, B => 
                           x_vector_91_port, ZN => mult_42_I10_n352);
   mult_42_I10_U386 : NAND2_X1 port map( A1 => mult_42_I10_n319, A2 => 
                           mult_42_I10_n402, ZN => mult_42_I10_n401);
   mult_42_I10_U385 : MUX2_X1 port map( A => mult_42_I10_n400, B => 
                           mult_42_I10_n401, S => B(90), Z => mult_42_I10_n396)
                           ;
   mult_42_I10_U384 : XOR2_X1 port map( A => x_vector_93_port, B => 
                           x_vector_92_port, Z => mult_42_I10_n399);
   mult_42_I10_U383 : NAND2_X1 port map( A1 => mult_42_I10_n352, A2 => 
                           mult_42_I10_n399, ZN => mult_42_I10_n351);
   mult_42_I10_U382 : NOR3_X1 port map( A1 => mult_42_I10_n352, A2 => B(90), A3
                           => mult_42_I10_n317, ZN => mult_42_I10_n398);
   mult_42_I10_U381 : AOI21_X1 port map( B1 => x_vector_93_port, B2 => 
                           mult_42_I10_n318, A => mult_42_I10_n398, ZN => 
                           mult_42_I10_n397);
   mult_42_I10_U380 : OAI222_X1 port map( A1 => mult_42_I10_n396, A2 => 
                           mult_42_I10_n311, B1 => mult_42_I10_n397, B2 => 
                           mult_42_I10_n396, C1 => mult_42_I10_n397, C2 => 
                           mult_42_I10_n311, ZN => mult_42_I10_n395);
   mult_42_I10_U379 : AOI222_X1 port map( A1 => mult_42_I10_n395, A2 => 
                           mult_42_I10_n88, B1 => mult_42_I10_n395, B2 => 
                           mult_42_I10_n89, C1 => mult_42_I10_n89, C2 => 
                           mult_42_I10_n88, ZN => mult_42_I10_n394);
   mult_42_I10_U378 : OAI222_X1 port map( A1 => mult_42_I10_n394, A2 => 
                           mult_42_I10_n308, B1 => mult_42_I10_n394, B2 => 
                           mult_42_I10_n309, C1 => mult_42_I10_n309, C2 => 
                           mult_42_I10_n308, ZN => mult_42_I10_n393);
   mult_42_I10_U377 : AOI222_X1 port map( A1 => mult_42_I10_n393, A2 => 
                           mult_42_I10_n80, B1 => mult_42_I10_n393, B2 => 
                           mult_42_I10_n83, C1 => mult_42_I10_n83, C2 => 
                           mult_42_I10_n80, ZN => mult_42_I10_n392);
   mult_42_I10_U376 : OAI222_X1 port map( A1 => mult_42_I10_n392, A2 => 
                           mult_42_I10_n305, B1 => mult_42_I10_n392, B2 => 
                           mult_42_I10_n307, C1 => mult_42_I10_n307, C2 => 
                           mult_42_I10_n305, ZN => mult_42_I10_n391);
   mult_42_I10_U375 : AOI222_X1 port map( A1 => mult_42_I10_n391, A2 => 
                           mult_42_I10_n68, B1 => mult_42_I10_n391, B2 => 
                           mult_42_I10_n73, C1 => mult_42_I10_n73, C2 => 
                           mult_42_I10_n68, ZN => mult_42_I10_n390);
   mult_42_I10_U374 : OAI222_X1 port map( A1 => mult_42_I10_n390, A2 => 
                           mult_42_I10_n296, B1 => mult_42_I10_n390, B2 => 
                           mult_42_I10_n304, C1 => mult_42_I10_n304, C2 => 
                           mult_42_I10_n296, ZN => mult_42_I10_n10);
   mult_42_I10_U373 : XOR2_X1 port map( A => x_vector_99_port, B => 
                           x_vector_98_port, Z => mult_42_I10_n389);
   mult_42_I10_U372 : NAND2_X1 port map( A1 => mult_42_I10_n338, A2 => 
                           mult_42_I10_n389, ZN => mult_42_I10_n337);
   mult_42_I10_U371 : OR3_X1 port map( A1 => mult_42_I10_n338, A2 => B(90), A3 
                           => mult_42_I10_n314, ZN => mult_42_I10_n388);
   mult_42_I10_U370 : OAI21_X1 port map( B1 => mult_42_I10_n314, B2 => 
                           mult_42_I10_n337, A => mult_42_I10_n388, ZN => 
                           mult_42_I10_n105);
   mult_42_I10_U369 : XOR2_X1 port map( A => x_vector_97_port, B => 
                           x_vector_96_port, Z => mult_42_I10_n387);
   mult_42_I10_U368 : NAND2_X1 port map( A1 => mult_42_I10_n327, A2 => 
                           mult_42_I10_n387, ZN => mult_42_I10_n326);
   mult_42_I10_U367 : OR3_X1 port map( A1 => mult_42_I10_n327, A2 => B(90), A3 
                           => mult_42_I10_n315, ZN => mult_42_I10_n386);
   mult_42_I10_U366 : OAI21_X1 port map( B1 => mult_42_I10_n315, B2 => 
                           mult_42_I10_n326, A => mult_42_I10_n386, ZN => 
                           mult_42_I10_n106);
   mult_42_I10_U365 : XOR2_X1 port map( A => x_vector_95_port, B => 
                           x_vector_94_port, Z => mult_42_I10_n385);
   mult_42_I10_U364 : NAND2_X1 port map( A1 => mult_42_I10_n332, A2 => 
                           mult_42_I10_n385, ZN => mult_42_I10_n331);
   mult_42_I10_U363 : OR3_X1 port map( A1 => mult_42_I10_n332, A2 => B(90), A3 
                           => mult_42_I10_n316, ZN => mult_42_I10_n384);
   mult_42_I10_U362 : OAI21_X1 port map( B1 => mult_42_I10_n316, B2 => 
                           mult_42_I10_n331, A => mult_42_I10_n384, ZN => 
                           mult_42_I10_n107);
   mult_42_I10_U361 : XOR2_X1 port map( A => B(99), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n339);
   mult_42_I10_U360 : OAI22_X1 port map( A1 => mult_42_I10_n339, A2 => 
                           mult_42_I10_n338, B1 => mult_42_I10_n337, B2 => 
                           mult_42_I10_n339, ZN => mult_42_I10_n383);
   mult_42_I10_U359 : XOR2_X1 port map( A => B(97), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n382);
   mult_42_I10_U358 : XOR2_X1 port map( A => B(98), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n336);
   mult_42_I10_U357 : OAI22_X1 port map( A1 => mult_42_I10_n382, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n336, ZN => mult_42_I10_n111);
   mult_42_I10_U356 : XOR2_X1 port map( A => B(96), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n381);
   mult_42_I10_U355 : OAI22_X1 port map( A1 => mult_42_I10_n381, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n382, ZN => mult_42_I10_n112);
   mult_42_I10_U354 : XOR2_X1 port map( A => B(95), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n380);
   mult_42_I10_U353 : OAI22_X1 port map( A1 => mult_42_I10_n380, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n381, ZN => mult_42_I10_n113);
   mult_42_I10_U352 : XOR2_X1 port map( A => B(94), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n379);
   mult_42_I10_U351 : OAI22_X1 port map( A1 => mult_42_I10_n379, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n380, ZN => mult_42_I10_n114);
   mult_42_I10_U350 : XOR2_X1 port map( A => B(93), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n378);
   mult_42_I10_U349 : OAI22_X1 port map( A1 => mult_42_I10_n378, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n379, ZN => mult_42_I10_n115);
   mult_42_I10_U348 : XOR2_X1 port map( A => B(92), B => mult_42_I10_n314, Z =>
                           mult_42_I10_n377);
   mult_42_I10_U347 : OAI22_X1 port map( A1 => mult_42_I10_n377, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n378, ZN => mult_42_I10_n116);
   mult_42_I10_U346 : XOR2_X1 port map( A => mult_42_I10_n312, B => 
                           x_vector_99_port, Z => mult_42_I10_n376);
   mult_42_I10_U345 : OAI22_X1 port map( A1 => mult_42_I10_n376, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n377, ZN => mult_42_I10_n117);
   mult_42_I10_U344 : XOR2_X1 port map( A => mult_42_I10_n314, B => B(90), Z =>
                           mult_42_I10_n375);
   mult_42_I10_U343 : OAI22_X1 port map( A1 => mult_42_I10_n375, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n376, ZN => mult_42_I10_n118);
   mult_42_I10_U342 : NOR2_X1 port map( A1 => mult_42_I10_n338, A2 => 
                           mult_42_I10_n313, ZN => mult_42_I10_n119);
   mult_42_I10_U341 : XOR2_X1 port map( A => B(99), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n335);
   mult_42_I10_U340 : OAI22_X1 port map( A1 => mult_42_I10_n335, A2 => 
                           mult_42_I10_n327, B1 => mult_42_I10_n326, B2 => 
                           mult_42_I10_n335, ZN => mult_42_I10_n374);
   mult_42_I10_U339 : XOR2_X1 port map( A => B(97), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n373);
   mult_42_I10_U338 : XOR2_X1 port map( A => B(98), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n334);
   mult_42_I10_U337 : OAI22_X1 port map( A1 => mult_42_I10_n373, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n334, ZN => mult_42_I10_n121);
   mult_42_I10_U336 : XOR2_X1 port map( A => B(96), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n372);
   mult_42_I10_U335 : OAI22_X1 port map( A1 => mult_42_I10_n372, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n373, ZN => mult_42_I10_n122);
   mult_42_I10_U334 : XOR2_X1 port map( A => B(95), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n371);
   mult_42_I10_U333 : OAI22_X1 port map( A1 => mult_42_I10_n371, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n372, ZN => mult_42_I10_n123);
   mult_42_I10_U332 : XOR2_X1 port map( A => B(94), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n328);
   mult_42_I10_U331 : OAI22_X1 port map( A1 => mult_42_I10_n328, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n371, ZN => mult_42_I10_n124);
   mult_42_I10_U330 : XOR2_X1 port map( A => B(92), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n370);
   mult_42_I10_U329 : XOR2_X1 port map( A => B(93), B => mult_42_I10_n315, Z =>
                           mult_42_I10_n325);
   mult_42_I10_U328 : OAI22_X1 port map( A1 => mult_42_I10_n370, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n325, ZN => mult_42_I10_n126);
   mult_42_I10_U327 : XOR2_X1 port map( A => mult_42_I10_n312, B => 
                           x_vector_97_port, Z => mult_42_I10_n369);
   mult_42_I10_U326 : OAI22_X1 port map( A1 => mult_42_I10_n369, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n370, ZN => mult_42_I10_n127);
   mult_42_I10_U325 : XOR2_X1 port map( A => mult_42_I10_n313, B => 
                           x_vector_97_port, Z => mult_42_I10_n368);
   mult_42_I10_U324 : OAI22_X1 port map( A1 => mult_42_I10_n368, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n369, ZN => mult_42_I10_n128);
   mult_42_I10_U323 : NOR2_X1 port map( A1 => mult_42_I10_n327, A2 => 
                           mult_42_I10_n313, ZN => mult_42_I10_n129);
   mult_42_I10_U322 : XOR2_X1 port map( A => B(99), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n333);
   mult_42_I10_U321 : OAI22_X1 port map( A1 => mult_42_I10_n333, A2 => 
                           mult_42_I10_n332, B1 => mult_42_I10_n331, B2 => 
                           mult_42_I10_n333, ZN => mult_42_I10_n367);
   mult_42_I10_U320 : XOR2_X1 port map( A => B(97), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n366);
   mult_42_I10_U319 : XOR2_X1 port map( A => B(98), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n330);
   mult_42_I10_U318 : OAI22_X1 port map( A1 => mult_42_I10_n366, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n330, ZN => mult_42_I10_n131);
   mult_42_I10_U317 : XOR2_X1 port map( A => B(96), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n365);
   mult_42_I10_U316 : OAI22_X1 port map( A1 => mult_42_I10_n365, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n366, ZN => mult_42_I10_n132);
   mult_42_I10_U315 : XOR2_X1 port map( A => B(95), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n364);
   mult_42_I10_U314 : OAI22_X1 port map( A1 => mult_42_I10_n364, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n365, ZN => mult_42_I10_n133);
   mult_42_I10_U313 : XOR2_X1 port map( A => B(94), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n363);
   mult_42_I10_U312 : OAI22_X1 port map( A1 => mult_42_I10_n363, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n364, ZN => mult_42_I10_n134);
   mult_42_I10_U311 : XOR2_X1 port map( A => B(93), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n362);
   mult_42_I10_U310 : OAI22_X1 port map( A1 => mult_42_I10_n362, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n363, ZN => mult_42_I10_n135);
   mult_42_I10_U309 : XOR2_X1 port map( A => B(92), B => mult_42_I10_n316, Z =>
                           mult_42_I10_n361);
   mult_42_I10_U308 : OAI22_X1 port map( A1 => mult_42_I10_n361, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n362, ZN => mult_42_I10_n136);
   mult_42_I10_U307 : XOR2_X1 port map( A => mult_42_I10_n312, B => 
                           x_vector_95_port, Z => mult_42_I10_n360);
   mult_42_I10_U306 : OAI22_X1 port map( A1 => mult_42_I10_n360, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n361, ZN => mult_42_I10_n137);
   mult_42_I10_U305 : XOR2_X1 port map( A => mult_42_I10_n313, B => 
                           x_vector_95_port, Z => mult_42_I10_n359);
   mult_42_I10_U304 : OAI22_X1 port map( A1 => mult_42_I10_n359, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n360, ZN => mult_42_I10_n138);
   mult_42_I10_U303 : NOR2_X1 port map( A1 => mult_42_I10_n332, A2 => 
                           mult_42_I10_n313, ZN => mult_42_I10_n139);
   mult_42_I10_U302 : XOR2_X1 port map( A => B(99), B => x_vector_93_port, Z =>
                           mult_42_I10_n329);
   mult_42_I10_U301 : AOI22_X1 port map( A1 => mult_42_I10_n329, A2 => 
                           mult_42_I10_n319, B1 => mult_42_I10_n318, B2 => 
                           mult_42_I10_n329, ZN => mult_42_I10_n140);
   mult_42_I10_U300 : XOR2_X1 port map( A => B(96), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n358);
   mult_42_I10_U299 : XOR2_X1 port map( A => B(97), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n324);
   mult_42_I10_U298 : OAI22_X1 port map( A1 => mult_42_I10_n358, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n324, ZN => mult_42_I10_n142);
   mult_42_I10_U297 : XOR2_X1 port map( A => B(95), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n357);
   mult_42_I10_U296 : OAI22_X1 port map( A1 => mult_42_I10_n357, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n358, ZN => mult_42_I10_n143);
   mult_42_I10_U295 : XOR2_X1 port map( A => B(94), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n356);
   mult_42_I10_U294 : OAI22_X1 port map( A1 => mult_42_I10_n356, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n357, ZN => mult_42_I10_n144);
   mult_42_I10_U293 : XOR2_X1 port map( A => B(93), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n355);
   mult_42_I10_U292 : OAI22_X1 port map( A1 => mult_42_I10_n355, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n356, ZN => mult_42_I10_n145);
   mult_42_I10_U291 : XOR2_X1 port map( A => B(92), B => mult_42_I10_n317, Z =>
                           mult_42_I10_n354);
   mult_42_I10_U290 : OAI22_X1 port map( A1 => mult_42_I10_n354, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n355, ZN => mult_42_I10_n146);
   mult_42_I10_U289 : XOR2_X1 port map( A => mult_42_I10_n312, B => 
                           x_vector_93_port, Z => mult_42_I10_n353);
   mult_42_I10_U288 : OAI22_X1 port map( A1 => mult_42_I10_n353, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n354, ZN => mult_42_I10_n147);
   mult_42_I10_U287 : XOR2_X1 port map( A => mult_42_I10_n313, B => 
                           x_vector_93_port, Z => mult_42_I10_n350);
   mult_42_I10_U286 : OAI22_X1 port map( A1 => mult_42_I10_n350, A2 => 
                           mult_42_I10_n351, B1 => mult_42_I10_n352, B2 => 
                           mult_42_I10_n353, ZN => mult_42_I10_n148);
   mult_42_I10_U285 : XNOR2_X1 port map( A => B(99), B => x_vector_91_port, ZN 
                           => mult_42_I10_n348);
   mult_42_I10_U284 : OAI22_X1 port map( A1 => mult_42_I10_n320, A2 => 
                           mult_42_I10_n348, B1 => mult_42_I10_n341, B2 => 
                           mult_42_I10_n348, ZN => mult_42_I10_n349);
   mult_42_I10_U283 : XNOR2_X1 port map( A => B(98), B => x_vector_91_port, ZN 
                           => mult_42_I10_n347);
   mult_42_I10_U282 : OAI22_X1 port map( A1 => mult_42_I10_n347, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n348, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n151);
   mult_42_I10_U281 : XNOR2_X1 port map( A => B(97), B => x_vector_91_port, ZN 
                           => mult_42_I10_n346);
   mult_42_I10_U280 : OAI22_X1 port map( A1 => mult_42_I10_n346, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n347, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n152);
   mult_42_I10_U279 : XNOR2_X1 port map( A => B(96), B => x_vector_91_port, ZN 
                           => mult_42_I10_n345);
   mult_42_I10_U278 : OAI22_X1 port map( A1 => mult_42_I10_n345, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n346, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n153);
   mult_42_I10_U277 : XNOR2_X1 port map( A => B(95), B => x_vector_91_port, ZN 
                           => mult_42_I10_n344);
   mult_42_I10_U276 : OAI22_X1 port map( A1 => mult_42_I10_n344, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n345, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n154);
   mult_42_I10_U275 : XNOR2_X1 port map( A => B(94), B => x_vector_91_port, ZN 
                           => mult_42_I10_n343);
   mult_42_I10_U274 : OAI22_X1 port map( A1 => mult_42_I10_n343, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n344, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n155);
   mult_42_I10_U273 : XNOR2_X1 port map( A => B(93), B => x_vector_91_port, ZN 
                           => mult_42_I10_n342);
   mult_42_I10_U272 : OAI22_X1 port map( A1 => mult_42_I10_n342, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n343, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n156);
   mult_42_I10_U271 : OAI22_X1 port map( A1 => mult_42_I10_n340, A2 => 
                           mult_42_I10_n341, B1 => mult_42_I10_n342, B2 => 
                           mult_42_I10_n320, ZN => mult_42_I10_n157);
   mult_42_I10_U270 : OAI22_X1 port map( A1 => mult_42_I10_n336, A2 => 
                           mult_42_I10_n337, B1 => mult_42_I10_n338, B2 => 
                           mult_42_I10_n339, ZN => mult_42_I10_n19);
   mult_42_I10_U269 : OAI22_X1 port map( A1 => mult_42_I10_n334, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n335, ZN => mult_42_I10_n25);
   mult_42_I10_U268 : OAI22_X1 port map( A1 => mult_42_I10_n330, A2 => 
                           mult_42_I10_n331, B1 => mult_42_I10_n332, B2 => 
                           mult_42_I10_n333, ZN => mult_42_I10_n35);
   mult_42_I10_U267 : XOR2_X1 port map( A => B(98), B => x_vector_93_port, Z =>
                           mult_42_I10_n323);
   mult_42_I10_U266 : AOI22_X1 port map( A1 => mult_42_I10_n323, A2 => 
                           mult_42_I10_n318, B1 => mult_42_I10_n319, B2 => 
                           mult_42_I10_n329, ZN => mult_42_I10_n50);
   mult_42_I10_U265 : OAI22_X1 port map( A1 => mult_42_I10_n325, A2 => 
                           mult_42_I10_n326, B1 => mult_42_I10_n327, B2 => 
                           mult_42_I10_n328, ZN => mult_42_I10_n321);
   mult_42_I10_U264 : AOI22_X1 port map( A1 => mult_42_I10_n306, A2 => 
                           mult_42_I10_n318, B1 => mult_42_I10_n319, B2 => 
                           mult_42_I10_n323, ZN => mult_42_I10_n322);
   mult_42_I10_U263 : NAND2_X1 port map( A1 => mult_42_I10_n310, A2 => 
                           mult_42_I10_n322, ZN => mult_42_I10_n57);
   mult_42_I10_U262 : XOR2_X1 port map( A => mult_42_I10_n321, B => 
                           mult_42_I10_n322, Z => mult_42_I10_n58);
   mult_42_I10_U261 : XNOR2_X2 port map( A => x_vector_98_port, B => 
                           x_vector_97_port, ZN => mult_42_I10_n338);
   mult_42_I10_U260 : XNOR2_X2 port map( A => x_vector_96_port, B => 
                           x_vector_95_port, ZN => mult_42_I10_n327);
   mult_42_I10_U259 : XNOR2_X2 port map( A => x_vector_94_port, B => 
                           x_vector_93_port, ZN => mult_42_I10_n332);
   mult_42_I10_U258 : INV_X1 port map( A => B(91), ZN => mult_42_I10_n312);
   mult_42_I10_U257 : INV_X1 port map( A => B(90), ZN => mult_42_I10_n313);
   mult_42_I10_U256 : INV_X1 port map( A => x_vector_93_port, ZN => 
                           mult_42_I10_n317);
   mult_42_I10_U255 : INV_X1 port map( A => x_vector_90_port, ZN => 
                           mult_42_I10_n320);
   mult_42_I10_U254 : INV_X1 port map( A => x_vector_97_port, ZN => 
                           mult_42_I10_n315);
   mult_42_I10_U253 : INV_X1 port map( A => x_vector_95_port, ZN => 
                           mult_42_I10_n316);
   mult_42_I10_U252 : INV_X1 port map( A => x_vector_99_port, ZN => 
                           mult_42_I10_n314);
   mult_42_I10_U251 : INV_X1 port map( A => mult_42_I10_n367, ZN => 
                           mult_42_I10_n298);
   mult_42_I10_U250 : INV_X1 port map( A => mult_42_I10_n374, ZN => 
                           mult_42_I10_n300);
   mult_42_I10_U249 : INV_X1 port map( A => mult_42_I10_n25, ZN => 
                           mult_42_I10_n301);
   mult_42_I10_U248 : INV_X1 port map( A => mult_42_I10_n35, ZN => 
                           mult_42_I10_n299);
   mult_42_I10_U247 : INV_X1 port map( A => mult_42_I10_n90, ZN => 
                           mult_42_I10_n311);
   mult_42_I10_U246 : INV_X1 port map( A => mult_42_I10_n50, ZN => 
                           mult_42_I10_n297);
   mult_42_I10_U245 : INV_X1 port map( A => mult_42_I10_n383, ZN => 
                           mult_42_I10_n302);
   mult_42_I10_U244 : INV_X1 port map( A => mult_42_I10_n349, ZN => 
                           mult_42_I10_n295);
   mult_42_I10_U243 : INV_X1 port map( A => mult_42_I10_n351, ZN => 
                           mult_42_I10_n318);
   mult_42_I10_U242 : INV_X1 port map( A => mult_42_I10_n352, ZN => 
                           mult_42_I10_n319);
   mult_42_I10_U241 : INV_X1 port map( A => mult_42_I10_n324, ZN => 
                           mult_42_I10_n306);
   mult_42_I10_U240 : INV_X1 port map( A => mult_42_I10_n84, ZN => 
                           mult_42_I10_n308);
   mult_42_I10_U239 : INV_X1 port map( A => mult_42_I10_n87, ZN => 
                           mult_42_I10_n309);
   mult_42_I10_U238 : INV_X1 port map( A => mult_42_I10_n19, ZN => 
                           mult_42_I10_n303);
   mult_42_I10_U237 : INV_X1 port map( A => mult_42_I10_n321, ZN => 
                           mult_42_I10_n310);
   mult_42_I10_U236 : INV_X1 port map( A => mult_42_I10_n1, ZN => N182_port);
   mult_42_I10_U235 : INV_X1 port map( A => mult_42_I10_n74, ZN => 
                           mult_42_I10_n305);
   mult_42_I10_U234 : INV_X1 port map( A => mult_42_I10_n79, ZN => 
                           mult_42_I10_n307);
   mult_42_I10_U233 : INV_X1 port map( A => mult_42_I10_n60, ZN => 
                           mult_42_I10_n296);
   mult_42_I10_U232 : INV_X1 port map( A => mult_42_I10_n67, ZN => 
                           mult_42_I10_n304);
   mult_42_I10_U56 : HA_X1 port map( A => mult_42_I10_n148, B => 
                           mult_42_I10_n157, CO => mult_42_I10_n89, S => 
                           mult_42_I10_n90);
   mult_42_I10_U55 : FA_X1 port map( A => mult_42_I10_n156, B => 
                           mult_42_I10_n139, CI => mult_42_I10_n147, CO => 
                           mult_42_I10_n87, S => mult_42_I10_n88);
   mult_42_I10_U54 : HA_X1 port map( A => mult_42_I10_n107, B => 
                           mult_42_I10_n138, CO => mult_42_I10_n85, S => 
                           mult_42_I10_n86);
   mult_42_I10_U53 : FA_X1 port map( A => mult_42_I10_n146, B => 
                           mult_42_I10_n155, CI => mult_42_I10_n86, CO => 
                           mult_42_I10_n83, S => mult_42_I10_n84);
   mult_42_I10_U52 : FA_X1 port map( A => mult_42_I10_n154, B => 
                           mult_42_I10_n129, CI => mult_42_I10_n145, CO => 
                           mult_42_I10_n81, S => mult_42_I10_n82);
   mult_42_I10_U51 : FA_X1 port map( A => mult_42_I10_n85, B => 
                           mult_42_I10_n137, CI => mult_42_I10_n82, CO => 
                           mult_42_I10_n79, S => mult_42_I10_n80);
   mult_42_I10_U50 : HA_X1 port map( A => mult_42_I10_n106, B => 
                           mult_42_I10_n128, CO => mult_42_I10_n77, S => 
                           mult_42_I10_n78);
   mult_42_I10_U49 : FA_X1 port map( A => mult_42_I10_n136, B => 
                           mult_42_I10_n153, CI => mult_42_I10_n144, CO => 
                           mult_42_I10_n75, S => mult_42_I10_n76);
   mult_42_I10_U48 : FA_X1 port map( A => mult_42_I10_n81, B => mult_42_I10_n78
                           , CI => mult_42_I10_n76, CO => mult_42_I10_n73, S =>
                           mult_42_I10_n74);
   mult_42_I10_U47 : FA_X1 port map( A => mult_42_I10_n135, B => 
                           mult_42_I10_n119, CI => mult_42_I10_n152, CO => 
                           mult_42_I10_n71, S => mult_42_I10_n72);
   mult_42_I10_U46 : FA_X1 port map( A => mult_42_I10_n127, B => 
                           mult_42_I10_n143, CI => mult_42_I10_n77, CO => 
                           mult_42_I10_n69, S => mult_42_I10_n70);
   mult_42_I10_U45 : FA_X1 port map( A => mult_42_I10_n72, B => mult_42_I10_n75
                           , CI => mult_42_I10_n70, CO => mult_42_I10_n67, S =>
                           mult_42_I10_n68);
   mult_42_I10_U44 : HA_X1 port map( A => mult_42_I10_n105, B => 
                           mult_42_I10_n118, CO => mult_42_I10_n65, S => 
                           mult_42_I10_n66);
   mult_42_I10_U43 : FA_X1 port map( A => mult_42_I10_n126, B => 
                           mult_42_I10_n134, CI => mult_42_I10_n142, CO => 
                           mult_42_I10_n63, S => mult_42_I10_n64);
   mult_42_I10_U42 : FA_X1 port map( A => mult_42_I10_n66, B => 
                           mult_42_I10_n151, CI => mult_42_I10_n71, CO => 
                           mult_42_I10_n61, S => mult_42_I10_n62);
   mult_42_I10_U41 : FA_X1 port map( A => mult_42_I10_n64, B => mult_42_I10_n69
                           , CI => mult_42_I10_n62, CO => mult_42_I10_n59, S =>
                           mult_42_I10_n60);
   mult_42_I10_U38 : FA_X1 port map( A => mult_42_I10_n133, B => 
                           mult_42_I10_n117, CI => mult_42_I10_n295, CO => 
                           mult_42_I10_n55, S => mult_42_I10_n56);
   mult_42_I10_U37 : FA_X1 port map( A => mult_42_I10_n58, B => mult_42_I10_n65
                           , CI => mult_42_I10_n63, CO => mult_42_I10_n53, S =>
                           mult_42_I10_n54);
   mult_42_I10_U36 : FA_X1 port map( A => mult_42_I10_n61, B => mult_42_I10_n56
                           , CI => mult_42_I10_n54, CO => mult_42_I10_n51, S =>
                           mult_42_I10_n52);
   mult_42_I10_U34 : FA_X1 port map( A => mult_42_I10_n124, B => 
                           mult_42_I10_n116, CI => mult_42_I10_n132, CO => 
                           mult_42_I10_n47, S => mult_42_I10_n48);
   mult_42_I10_U33 : FA_X1 port map( A => mult_42_I10_n57, B => mult_42_I10_n50
                           , CI => mult_42_I10_n55, CO => mult_42_I10_n45, S =>
                           mult_42_I10_n46);
   mult_42_I10_U32 : FA_X1 port map( A => mult_42_I10_n53, B => mult_42_I10_n48
                           , CI => mult_42_I10_n46, CO => mult_42_I10_n43, S =>
                           mult_42_I10_n44);
   mult_42_I10_U31 : FA_X1 port map( A => mult_42_I10_n123, B => 
                           mult_42_I10_n115, CI => mult_42_I10_n140, CO => 
                           mult_42_I10_n41, S => mult_42_I10_n42);
   mult_42_I10_U30 : FA_X1 port map( A => mult_42_I10_n297, B => 
                           mult_42_I10_n131, CI => mult_42_I10_n47, CO => 
                           mult_42_I10_n39, S => mult_42_I10_n40);
   mult_42_I10_U29 : FA_X1 port map( A => mult_42_I10_n45, B => mult_42_I10_n42
                           , CI => mult_42_I10_n40, CO => mult_42_I10_n37, S =>
                           mult_42_I10_n38);
   mult_42_I10_U27 : FA_X1 port map( A => mult_42_I10_n114, B => 
                           mult_42_I10_n122, CI => mult_42_I10_n299, CO => 
                           mult_42_I10_n33, S => mult_42_I10_n34);
   mult_42_I10_U26 : FA_X1 port map( A => mult_42_I10_n34, B => mult_42_I10_n41
                           , CI => mult_42_I10_n39, CO => mult_42_I10_n31, S =>
                           mult_42_I10_n32);
   mult_42_I10_U25 : FA_X1 port map( A => mult_42_I10_n121, B => 
                           mult_42_I10_n35, CI => mult_42_I10_n298, CO => 
                           mult_42_I10_n29, S => mult_42_I10_n30);
   mult_42_I10_U24 : FA_X1 port map( A => mult_42_I10_n33, B => 
                           mult_42_I10_n113, CI => mult_42_I10_n30, CO => 
                           mult_42_I10_n27, S => mult_42_I10_n28);
   mult_42_I10_U22 : FA_X1 port map( A => mult_42_I10_n301, B => 
                           mult_42_I10_n112, CI => mult_42_I10_n29, CO => 
                           mult_42_I10_n23, S => mult_42_I10_n24);
   mult_42_I10_U21 : FA_X1 port map( A => mult_42_I10_n111, B => 
                           mult_42_I10_n25, CI => mult_42_I10_n300, CO => 
                           mult_42_I10_n21, S => mult_42_I10_n22);
   mult_42_I10_U10 : FA_X1 port map( A => mult_42_I10_n52, B => mult_42_I10_n59
                           , CI => mult_42_I10_n10, CO => mult_42_I10_n9, S => 
                           N173_port);
   mult_42_I10_U9 : FA_X1 port map( A => mult_42_I10_n44, B => mult_42_I10_n51,
                           CI => mult_42_I10_n9, CO => mult_42_I10_n8, S => 
                           N174_port);
   mult_42_I10_U8 : FA_X1 port map( A => mult_42_I10_n38, B => mult_42_I10_n43,
                           CI => mult_42_I10_n8, CO => mult_42_I10_n7, S => 
                           N175_port);
   mult_42_I10_U7 : FA_X1 port map( A => mult_42_I10_n32, B => mult_42_I10_n37,
                           CI => mult_42_I10_n7, CO => mult_42_I10_n6, S => 
                           N176_port);
   mult_42_I10_U6 : FA_X1 port map( A => mult_42_I10_n28, B => mult_42_I10_n31,
                           CI => mult_42_I10_n6, CO => mult_42_I10_n5, S => 
                           N177_port);
   mult_42_I10_U5 : FA_X1 port map( A => mult_42_I10_n24, B => mult_42_I10_n27,
                           CI => mult_42_I10_n5, CO => mult_42_I10_n4, S => 
                           N178_port);
   mult_42_I10_U4 : FA_X1 port map( A => mult_42_I10_n23, B => mult_42_I10_n22,
                           CI => mult_42_I10_n4, CO => mult_42_I10_n3, S => 
                           N179_port);
   mult_42_I10_U3 : FA_X1 port map( A => mult_42_I10_n21, B => mult_42_I10_n303
                           , CI => mult_42_I10_n3, CO => mult_42_I10_n2, S => 
                           N180_port);
   mult_42_I10_U2 : FA_X1 port map( A => mult_42_I10_n302, B => mult_42_I10_n19
                           , CI => mult_42_I10_n2, CO => mult_42_I10_n1, S => 
                           N181_port);
   mult_42_I11_U391 : NAND2_X1 port map( A1 => x_vector_101_port, A2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n341);
   mult_42_I11_U390 : XNOR2_X1 port map( A => B(102), B => x_vector_101_port, 
                           ZN => mult_42_I11_n340);
   mult_42_I11_U389 : OAI22_X1 port map( A1 => B(101), A2 => mult_42_I11_n341, 
                           B1 => mult_42_I11_n340, B2 => mult_42_I11_n320, ZN 
                           => mult_42_I11_n402);
   mult_42_I11_U388 : NAND3_X1 port map( A1 => mult_42_I11_n402, A2 => 
                           mult_42_I11_n312, A3 => x_vector_101_port, ZN => 
                           mult_42_I11_n400);
   mult_42_I11_U387 : XNOR2_X1 port map( A => x_vector_102_port, B => 
                           x_vector_101_port, ZN => mult_42_I11_n352);
   mult_42_I11_U386 : NAND2_X1 port map( A1 => mult_42_I11_n319, A2 => 
                           mult_42_I11_n402, ZN => mult_42_I11_n401);
   mult_42_I11_U385 : MUX2_X1 port map( A => mult_42_I11_n400, B => 
                           mult_42_I11_n401, S => B(100), Z => mult_42_I11_n396
                           );
   mult_42_I11_U384 : XOR2_X1 port map( A => x_vector_103_port, B => 
                           x_vector_102_port, Z => mult_42_I11_n399);
   mult_42_I11_U383 : NAND2_X1 port map( A1 => mult_42_I11_n352, A2 => 
                           mult_42_I11_n399, ZN => mult_42_I11_n351);
   mult_42_I11_U382 : NOR3_X1 port map( A1 => mult_42_I11_n352, A2 => B(100), 
                           A3 => mult_42_I11_n317, ZN => mult_42_I11_n398);
   mult_42_I11_U381 : AOI21_X1 port map( B1 => x_vector_103_port, B2 => 
                           mult_42_I11_n318, A => mult_42_I11_n398, ZN => 
                           mult_42_I11_n397);
   mult_42_I11_U380 : OAI222_X1 port map( A1 => mult_42_I11_n396, A2 => 
                           mult_42_I11_n311, B1 => mult_42_I11_n397, B2 => 
                           mult_42_I11_n396, C1 => mult_42_I11_n397, C2 => 
                           mult_42_I11_n311, ZN => mult_42_I11_n395);
   mult_42_I11_U379 : AOI222_X1 port map( A1 => mult_42_I11_n395, A2 => 
                           mult_42_I11_n88, B1 => mult_42_I11_n395, B2 => 
                           mult_42_I11_n89, C1 => mult_42_I11_n89, C2 => 
                           mult_42_I11_n88, ZN => mult_42_I11_n394);
   mult_42_I11_U378 : OAI222_X1 port map( A1 => mult_42_I11_n394, A2 => 
                           mult_42_I11_n308, B1 => mult_42_I11_n394, B2 => 
                           mult_42_I11_n309, C1 => mult_42_I11_n309, C2 => 
                           mult_42_I11_n308, ZN => mult_42_I11_n393);
   mult_42_I11_U377 : AOI222_X1 port map( A1 => mult_42_I11_n393, A2 => 
                           mult_42_I11_n80, B1 => mult_42_I11_n393, B2 => 
                           mult_42_I11_n83, C1 => mult_42_I11_n83, C2 => 
                           mult_42_I11_n80, ZN => mult_42_I11_n392);
   mult_42_I11_U376 : OAI222_X1 port map( A1 => mult_42_I11_n392, A2 => 
                           mult_42_I11_n305, B1 => mult_42_I11_n392, B2 => 
                           mult_42_I11_n307, C1 => mult_42_I11_n307, C2 => 
                           mult_42_I11_n305, ZN => mult_42_I11_n391);
   mult_42_I11_U375 : AOI222_X1 port map( A1 => mult_42_I11_n391, A2 => 
                           mult_42_I11_n68, B1 => mult_42_I11_n391, B2 => 
                           mult_42_I11_n73, C1 => mult_42_I11_n73, C2 => 
                           mult_42_I11_n68, ZN => mult_42_I11_n390);
   mult_42_I11_U374 : OAI222_X1 port map( A1 => mult_42_I11_n390, A2 => 
                           mult_42_I11_n296, B1 => mult_42_I11_n390, B2 => 
                           mult_42_I11_n304, C1 => mult_42_I11_n304, C2 => 
                           mult_42_I11_n296, ZN => mult_42_I11_n10);
   mult_42_I11_U373 : XOR2_X1 port map( A => x_vector_109_port, B => 
                           x_vector_108_port, Z => mult_42_I11_n389);
   mult_42_I11_U372 : NAND2_X1 port map( A1 => mult_42_I11_n338, A2 => 
                           mult_42_I11_n389, ZN => mult_42_I11_n337);
   mult_42_I11_U371 : OR3_X1 port map( A1 => mult_42_I11_n338, A2 => B(100), A3
                           => mult_42_I11_n314, ZN => mult_42_I11_n388);
   mult_42_I11_U370 : OAI21_X1 port map( B1 => mult_42_I11_n314, B2 => 
                           mult_42_I11_n337, A => mult_42_I11_n388, ZN => 
                           mult_42_I11_n105);
   mult_42_I11_U369 : XOR2_X1 port map( A => x_vector_107_port, B => 
                           x_vector_106_port, Z => mult_42_I11_n387);
   mult_42_I11_U368 : NAND2_X1 port map( A1 => mult_42_I11_n327, A2 => 
                           mult_42_I11_n387, ZN => mult_42_I11_n326);
   mult_42_I11_U367 : OR3_X1 port map( A1 => mult_42_I11_n327, A2 => B(100), A3
                           => mult_42_I11_n315, ZN => mult_42_I11_n386);
   mult_42_I11_U366 : OAI21_X1 port map( B1 => mult_42_I11_n315, B2 => 
                           mult_42_I11_n326, A => mult_42_I11_n386, ZN => 
                           mult_42_I11_n106);
   mult_42_I11_U365 : XOR2_X1 port map( A => x_vector_105_port, B => 
                           x_vector_104_port, Z => mult_42_I11_n385);
   mult_42_I11_U364 : NAND2_X1 port map( A1 => mult_42_I11_n332, A2 => 
                           mult_42_I11_n385, ZN => mult_42_I11_n331);
   mult_42_I11_U363 : OR3_X1 port map( A1 => mult_42_I11_n332, A2 => B(100), A3
                           => mult_42_I11_n316, ZN => mult_42_I11_n384);
   mult_42_I11_U362 : OAI21_X1 port map( B1 => mult_42_I11_n316, B2 => 
                           mult_42_I11_n331, A => mult_42_I11_n384, ZN => 
                           mult_42_I11_n107);
   mult_42_I11_U361 : XOR2_X1 port map( A => B(109), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n339);
   mult_42_I11_U360 : OAI22_X1 port map( A1 => mult_42_I11_n339, A2 => 
                           mult_42_I11_n338, B1 => mult_42_I11_n337, B2 => 
                           mult_42_I11_n339, ZN => mult_42_I11_n383);
   mult_42_I11_U359 : XOR2_X1 port map( A => B(107), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n382);
   mult_42_I11_U358 : XOR2_X1 port map( A => B(108), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n336);
   mult_42_I11_U357 : OAI22_X1 port map( A1 => mult_42_I11_n382, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n336, ZN => mult_42_I11_n111);
   mult_42_I11_U356 : XOR2_X1 port map( A => B(106), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n381);
   mult_42_I11_U355 : OAI22_X1 port map( A1 => mult_42_I11_n381, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n382, ZN => mult_42_I11_n112);
   mult_42_I11_U354 : XOR2_X1 port map( A => B(105), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n380);
   mult_42_I11_U353 : OAI22_X1 port map( A1 => mult_42_I11_n380, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n381, ZN => mult_42_I11_n113);
   mult_42_I11_U352 : XOR2_X1 port map( A => B(104), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n379);
   mult_42_I11_U351 : OAI22_X1 port map( A1 => mult_42_I11_n379, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n380, ZN => mult_42_I11_n114);
   mult_42_I11_U350 : XOR2_X1 port map( A => B(103), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n378);
   mult_42_I11_U349 : OAI22_X1 port map( A1 => mult_42_I11_n378, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n379, ZN => mult_42_I11_n115);
   mult_42_I11_U348 : XOR2_X1 port map( A => B(102), B => mult_42_I11_n314, Z 
                           => mult_42_I11_n377);
   mult_42_I11_U347 : OAI22_X1 port map( A1 => mult_42_I11_n377, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n378, ZN => mult_42_I11_n116);
   mult_42_I11_U346 : XOR2_X1 port map( A => mult_42_I11_n312, B => 
                           x_vector_109_port, Z => mult_42_I11_n376);
   mult_42_I11_U345 : OAI22_X1 port map( A1 => mult_42_I11_n376, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n377, ZN => mult_42_I11_n117);
   mult_42_I11_U344 : XOR2_X1 port map( A => mult_42_I11_n314, B => B(100), Z 
                           => mult_42_I11_n375);
   mult_42_I11_U343 : OAI22_X1 port map( A1 => mult_42_I11_n375, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n376, ZN => mult_42_I11_n118);
   mult_42_I11_U342 : NOR2_X1 port map( A1 => mult_42_I11_n338, A2 => 
                           mult_42_I11_n313, ZN => mult_42_I11_n119);
   mult_42_I11_U341 : XOR2_X1 port map( A => B(109), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n335);
   mult_42_I11_U340 : OAI22_X1 port map( A1 => mult_42_I11_n335, A2 => 
                           mult_42_I11_n327, B1 => mult_42_I11_n326, B2 => 
                           mult_42_I11_n335, ZN => mult_42_I11_n374);
   mult_42_I11_U339 : XOR2_X1 port map( A => B(107), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n373);
   mult_42_I11_U338 : XOR2_X1 port map( A => B(108), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n334);
   mult_42_I11_U337 : OAI22_X1 port map( A1 => mult_42_I11_n373, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n334, ZN => mult_42_I11_n121);
   mult_42_I11_U336 : XOR2_X1 port map( A => B(106), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n372);
   mult_42_I11_U335 : OAI22_X1 port map( A1 => mult_42_I11_n372, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n373, ZN => mult_42_I11_n122);
   mult_42_I11_U334 : XOR2_X1 port map( A => B(105), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n371);
   mult_42_I11_U333 : OAI22_X1 port map( A1 => mult_42_I11_n371, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n372, ZN => mult_42_I11_n123);
   mult_42_I11_U332 : XOR2_X1 port map( A => B(104), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n328);
   mult_42_I11_U331 : OAI22_X1 port map( A1 => mult_42_I11_n328, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n371, ZN => mult_42_I11_n124);
   mult_42_I11_U330 : XOR2_X1 port map( A => B(102), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n370);
   mult_42_I11_U329 : XOR2_X1 port map( A => B(103), B => mult_42_I11_n315, Z 
                           => mult_42_I11_n325);
   mult_42_I11_U328 : OAI22_X1 port map( A1 => mult_42_I11_n370, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n325, ZN => mult_42_I11_n126);
   mult_42_I11_U327 : XOR2_X1 port map( A => mult_42_I11_n312, B => 
                           x_vector_107_port, Z => mult_42_I11_n369);
   mult_42_I11_U326 : OAI22_X1 port map( A1 => mult_42_I11_n369, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n370, ZN => mult_42_I11_n127);
   mult_42_I11_U325 : XOR2_X1 port map( A => mult_42_I11_n313, B => 
                           x_vector_107_port, Z => mult_42_I11_n368);
   mult_42_I11_U324 : OAI22_X1 port map( A1 => mult_42_I11_n368, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n369, ZN => mult_42_I11_n128);
   mult_42_I11_U323 : NOR2_X1 port map( A1 => mult_42_I11_n327, A2 => 
                           mult_42_I11_n313, ZN => mult_42_I11_n129);
   mult_42_I11_U322 : XOR2_X1 port map( A => B(109), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n333);
   mult_42_I11_U321 : OAI22_X1 port map( A1 => mult_42_I11_n333, A2 => 
                           mult_42_I11_n332, B1 => mult_42_I11_n331, B2 => 
                           mult_42_I11_n333, ZN => mult_42_I11_n367);
   mult_42_I11_U320 : XOR2_X1 port map( A => B(107), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n366);
   mult_42_I11_U319 : XOR2_X1 port map( A => B(108), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n330);
   mult_42_I11_U318 : OAI22_X1 port map( A1 => mult_42_I11_n366, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n330, ZN => mult_42_I11_n131);
   mult_42_I11_U317 : XOR2_X1 port map( A => B(106), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n365);
   mult_42_I11_U316 : OAI22_X1 port map( A1 => mult_42_I11_n365, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n366, ZN => mult_42_I11_n132);
   mult_42_I11_U315 : XOR2_X1 port map( A => B(105), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n364);
   mult_42_I11_U314 : OAI22_X1 port map( A1 => mult_42_I11_n364, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n365, ZN => mult_42_I11_n133);
   mult_42_I11_U313 : XOR2_X1 port map( A => B(104), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n363);
   mult_42_I11_U312 : OAI22_X1 port map( A1 => mult_42_I11_n363, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n364, ZN => mult_42_I11_n134);
   mult_42_I11_U311 : XOR2_X1 port map( A => B(103), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n362);
   mult_42_I11_U310 : OAI22_X1 port map( A1 => mult_42_I11_n362, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n363, ZN => mult_42_I11_n135);
   mult_42_I11_U309 : XOR2_X1 port map( A => B(102), B => mult_42_I11_n316, Z 
                           => mult_42_I11_n361);
   mult_42_I11_U308 : OAI22_X1 port map( A1 => mult_42_I11_n361, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n362, ZN => mult_42_I11_n136);
   mult_42_I11_U307 : XOR2_X1 port map( A => mult_42_I11_n312, B => 
                           x_vector_105_port, Z => mult_42_I11_n360);
   mult_42_I11_U306 : OAI22_X1 port map( A1 => mult_42_I11_n360, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n361, ZN => mult_42_I11_n137);
   mult_42_I11_U305 : XOR2_X1 port map( A => mult_42_I11_n313, B => 
                           x_vector_105_port, Z => mult_42_I11_n359);
   mult_42_I11_U304 : OAI22_X1 port map( A1 => mult_42_I11_n359, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n360, ZN => mult_42_I11_n138);
   mult_42_I11_U303 : NOR2_X1 port map( A1 => mult_42_I11_n332, A2 => 
                           mult_42_I11_n313, ZN => mult_42_I11_n139);
   mult_42_I11_U302 : XOR2_X1 port map( A => B(109), B => x_vector_103_port, Z 
                           => mult_42_I11_n329);
   mult_42_I11_U301 : AOI22_X1 port map( A1 => mult_42_I11_n329, A2 => 
                           mult_42_I11_n319, B1 => mult_42_I11_n318, B2 => 
                           mult_42_I11_n329, ZN => mult_42_I11_n140);
   mult_42_I11_U300 : XOR2_X1 port map( A => B(106), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n358);
   mult_42_I11_U299 : XOR2_X1 port map( A => B(107), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n324);
   mult_42_I11_U298 : OAI22_X1 port map( A1 => mult_42_I11_n358, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n324, ZN => mult_42_I11_n142);
   mult_42_I11_U297 : XOR2_X1 port map( A => B(105), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n357);
   mult_42_I11_U296 : OAI22_X1 port map( A1 => mult_42_I11_n357, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n358, ZN => mult_42_I11_n143);
   mult_42_I11_U295 : XOR2_X1 port map( A => B(104), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n356);
   mult_42_I11_U294 : OAI22_X1 port map( A1 => mult_42_I11_n356, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n357, ZN => mult_42_I11_n144);
   mult_42_I11_U293 : XOR2_X1 port map( A => B(103), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n355);
   mult_42_I11_U292 : OAI22_X1 port map( A1 => mult_42_I11_n355, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n356, ZN => mult_42_I11_n145);
   mult_42_I11_U291 : XOR2_X1 port map( A => B(102), B => mult_42_I11_n317, Z 
                           => mult_42_I11_n354);
   mult_42_I11_U290 : OAI22_X1 port map( A1 => mult_42_I11_n354, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n355, ZN => mult_42_I11_n146);
   mult_42_I11_U289 : XOR2_X1 port map( A => mult_42_I11_n312, B => 
                           x_vector_103_port, Z => mult_42_I11_n353);
   mult_42_I11_U288 : OAI22_X1 port map( A1 => mult_42_I11_n353, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n354, ZN => mult_42_I11_n147);
   mult_42_I11_U287 : XOR2_X1 port map( A => mult_42_I11_n313, B => 
                           x_vector_103_port, Z => mult_42_I11_n350);
   mult_42_I11_U286 : OAI22_X1 port map( A1 => mult_42_I11_n350, A2 => 
                           mult_42_I11_n351, B1 => mult_42_I11_n352, B2 => 
                           mult_42_I11_n353, ZN => mult_42_I11_n148);
   mult_42_I11_U285 : XNOR2_X1 port map( A => B(109), B => x_vector_101_port, 
                           ZN => mult_42_I11_n348);
   mult_42_I11_U284 : OAI22_X1 port map( A1 => mult_42_I11_n320, A2 => 
                           mult_42_I11_n348, B1 => mult_42_I11_n341, B2 => 
                           mult_42_I11_n348, ZN => mult_42_I11_n349);
   mult_42_I11_U283 : XNOR2_X1 port map( A => B(108), B => x_vector_101_port, 
                           ZN => mult_42_I11_n347);
   mult_42_I11_U282 : OAI22_X1 port map( A1 => mult_42_I11_n347, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n348, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n151);
   mult_42_I11_U281 : XNOR2_X1 port map( A => B(107), B => x_vector_101_port, 
                           ZN => mult_42_I11_n346);
   mult_42_I11_U280 : OAI22_X1 port map( A1 => mult_42_I11_n346, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n347, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n152);
   mult_42_I11_U279 : XNOR2_X1 port map( A => B(106), B => x_vector_101_port, 
                           ZN => mult_42_I11_n345);
   mult_42_I11_U278 : OAI22_X1 port map( A1 => mult_42_I11_n345, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n346, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n153);
   mult_42_I11_U277 : XNOR2_X1 port map( A => B(105), B => x_vector_101_port, 
                           ZN => mult_42_I11_n344);
   mult_42_I11_U276 : OAI22_X1 port map( A1 => mult_42_I11_n344, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n345, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n154);
   mult_42_I11_U275 : XNOR2_X1 port map( A => B(104), B => x_vector_101_port, 
                           ZN => mult_42_I11_n343);
   mult_42_I11_U274 : OAI22_X1 port map( A1 => mult_42_I11_n343, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n344, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n155);
   mult_42_I11_U273 : XNOR2_X1 port map( A => B(103), B => x_vector_101_port, 
                           ZN => mult_42_I11_n342);
   mult_42_I11_U272 : OAI22_X1 port map( A1 => mult_42_I11_n342, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n343, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n156);
   mult_42_I11_U271 : OAI22_X1 port map( A1 => mult_42_I11_n340, A2 => 
                           mult_42_I11_n341, B1 => mult_42_I11_n342, B2 => 
                           mult_42_I11_n320, ZN => mult_42_I11_n157);
   mult_42_I11_U270 : OAI22_X1 port map( A1 => mult_42_I11_n336, A2 => 
                           mult_42_I11_n337, B1 => mult_42_I11_n338, B2 => 
                           mult_42_I11_n339, ZN => mult_42_I11_n19);
   mult_42_I11_U269 : OAI22_X1 port map( A1 => mult_42_I11_n334, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n335, ZN => mult_42_I11_n25);
   mult_42_I11_U268 : OAI22_X1 port map( A1 => mult_42_I11_n330, A2 => 
                           mult_42_I11_n331, B1 => mult_42_I11_n332, B2 => 
                           mult_42_I11_n333, ZN => mult_42_I11_n35);
   mult_42_I11_U267 : XOR2_X1 port map( A => B(108), B => x_vector_103_port, Z 
                           => mult_42_I11_n323);
   mult_42_I11_U266 : AOI22_X1 port map( A1 => mult_42_I11_n323, A2 => 
                           mult_42_I11_n318, B1 => mult_42_I11_n319, B2 => 
                           mult_42_I11_n329, ZN => mult_42_I11_n50);
   mult_42_I11_U265 : OAI22_X1 port map( A1 => mult_42_I11_n325, A2 => 
                           mult_42_I11_n326, B1 => mult_42_I11_n327, B2 => 
                           mult_42_I11_n328, ZN => mult_42_I11_n321);
   mult_42_I11_U264 : AOI22_X1 port map( A1 => mult_42_I11_n306, A2 => 
                           mult_42_I11_n318, B1 => mult_42_I11_n319, B2 => 
                           mult_42_I11_n323, ZN => mult_42_I11_n322);
   mult_42_I11_U263 : NAND2_X1 port map( A1 => mult_42_I11_n310, A2 => 
                           mult_42_I11_n322, ZN => mult_42_I11_n57);
   mult_42_I11_U262 : XOR2_X1 port map( A => mult_42_I11_n321, B => 
                           mult_42_I11_n322, Z => mult_42_I11_n58);
   mult_42_I11_U261 : XNOR2_X2 port map( A => x_vector_108_port, B => 
                           x_vector_107_port, ZN => mult_42_I11_n338);
   mult_42_I11_U260 : XNOR2_X2 port map( A => x_vector_106_port, B => 
                           x_vector_105_port, ZN => mult_42_I11_n327);
   mult_42_I11_U259 : XNOR2_X2 port map( A => x_vector_104_port, B => 
                           x_vector_103_port, ZN => mult_42_I11_n332);
   mult_42_I11_U258 : INV_X1 port map( A => B(101), ZN => mult_42_I11_n312);
   mult_42_I11_U257 : INV_X1 port map( A => B(100), ZN => mult_42_I11_n313);
   mult_42_I11_U256 : INV_X1 port map( A => x_vector_103_port, ZN => 
                           mult_42_I11_n317);
   mult_42_I11_U255 : INV_X1 port map( A => x_vector_100_port, ZN => 
                           mult_42_I11_n320);
   mult_42_I11_U254 : INV_X1 port map( A => x_vector_107_port, ZN => 
                           mult_42_I11_n315);
   mult_42_I11_U253 : INV_X1 port map( A => x_vector_105_port, ZN => 
                           mult_42_I11_n316);
   mult_42_I11_U252 : INV_X1 port map( A => x_vector_109_port, ZN => 
                           mult_42_I11_n314);
   mult_42_I11_U251 : INV_X1 port map( A => mult_42_I11_n374, ZN => 
                           mult_42_I11_n300);
   mult_42_I11_U250 : INV_X1 port map( A => mult_42_I11_n25, ZN => 
                           mult_42_I11_n301);
   mult_42_I11_U249 : INV_X1 port map( A => mult_42_I11_n90, ZN => 
                           mult_42_I11_n311);
   mult_42_I11_U248 : INV_X1 port map( A => mult_42_I11_n50, ZN => 
                           mult_42_I11_n297);
   mult_42_I11_U247 : INV_X1 port map( A => mult_42_I11_n367, ZN => 
                           mult_42_I11_n298);
   mult_42_I11_U246 : INV_X1 port map( A => mult_42_I11_n383, ZN => 
                           mult_42_I11_n302);
   mult_42_I11_U245 : INV_X1 port map( A => mult_42_I11_n349, ZN => 
                           mult_42_I11_n295);
   mult_42_I11_U244 : INV_X1 port map( A => mult_42_I11_n35, ZN => 
                           mult_42_I11_n299);
   mult_42_I11_U243 : INV_X1 port map( A => mult_42_I11_n351, ZN => 
                           mult_42_I11_n318);
   mult_42_I11_U242 : INV_X1 port map( A => mult_42_I11_n352, ZN => 
                           mult_42_I11_n319);
   mult_42_I11_U241 : INV_X1 port map( A => mult_42_I11_n324, ZN => 
                           mult_42_I11_n306);
   mult_42_I11_U240 : INV_X1 port map( A => mult_42_I11_n84, ZN => 
                           mult_42_I11_n308);
   mult_42_I11_U239 : INV_X1 port map( A => mult_42_I11_n87, ZN => 
                           mult_42_I11_n309);
   mult_42_I11_U238 : INV_X1 port map( A => mult_42_I11_n19, ZN => 
                           mult_42_I11_n303);
   mult_42_I11_U237 : INV_X1 port map( A => mult_42_I11_n321, ZN => 
                           mult_42_I11_n310);
   mult_42_I11_U236 : INV_X1 port map( A => mult_42_I11_n1, ZN => N202_port);
   mult_42_I11_U235 : INV_X1 port map( A => mult_42_I11_n74, ZN => 
                           mult_42_I11_n305);
   mult_42_I11_U234 : INV_X1 port map( A => mult_42_I11_n79, ZN => 
                           mult_42_I11_n307);
   mult_42_I11_U233 : INV_X1 port map( A => mult_42_I11_n60, ZN => 
                           mult_42_I11_n296);
   mult_42_I11_U232 : INV_X1 port map( A => mult_42_I11_n67, ZN => 
                           mult_42_I11_n304);
   mult_42_I11_U56 : HA_X1 port map( A => mult_42_I11_n148, B => 
                           mult_42_I11_n157, CO => mult_42_I11_n89, S => 
                           mult_42_I11_n90);
   mult_42_I11_U55 : FA_X1 port map( A => mult_42_I11_n156, B => 
                           mult_42_I11_n139, CI => mult_42_I11_n147, CO => 
                           mult_42_I11_n87, S => mult_42_I11_n88);
   mult_42_I11_U54 : HA_X1 port map( A => mult_42_I11_n107, B => 
                           mult_42_I11_n138, CO => mult_42_I11_n85, S => 
                           mult_42_I11_n86);
   mult_42_I11_U53 : FA_X1 port map( A => mult_42_I11_n146, B => 
                           mult_42_I11_n155, CI => mult_42_I11_n86, CO => 
                           mult_42_I11_n83, S => mult_42_I11_n84);
   mult_42_I11_U52 : FA_X1 port map( A => mult_42_I11_n154, B => 
                           mult_42_I11_n129, CI => mult_42_I11_n145, CO => 
                           mult_42_I11_n81, S => mult_42_I11_n82);
   mult_42_I11_U51 : FA_X1 port map( A => mult_42_I11_n85, B => 
                           mult_42_I11_n137, CI => mult_42_I11_n82, CO => 
                           mult_42_I11_n79, S => mult_42_I11_n80);
   mult_42_I11_U50 : HA_X1 port map( A => mult_42_I11_n106, B => 
                           mult_42_I11_n128, CO => mult_42_I11_n77, S => 
                           mult_42_I11_n78);
   mult_42_I11_U49 : FA_X1 port map( A => mult_42_I11_n136, B => 
                           mult_42_I11_n153, CI => mult_42_I11_n144, CO => 
                           mult_42_I11_n75, S => mult_42_I11_n76);
   mult_42_I11_U48 : FA_X1 port map( A => mult_42_I11_n81, B => mult_42_I11_n78
                           , CI => mult_42_I11_n76, CO => mult_42_I11_n73, S =>
                           mult_42_I11_n74);
   mult_42_I11_U47 : FA_X1 port map( A => mult_42_I11_n135, B => 
                           mult_42_I11_n119, CI => mult_42_I11_n152, CO => 
                           mult_42_I11_n71, S => mult_42_I11_n72);
   mult_42_I11_U46 : FA_X1 port map( A => mult_42_I11_n127, B => 
                           mult_42_I11_n143, CI => mult_42_I11_n77, CO => 
                           mult_42_I11_n69, S => mult_42_I11_n70);
   mult_42_I11_U45 : FA_X1 port map( A => mult_42_I11_n72, B => mult_42_I11_n75
                           , CI => mult_42_I11_n70, CO => mult_42_I11_n67, S =>
                           mult_42_I11_n68);
   mult_42_I11_U44 : HA_X1 port map( A => mult_42_I11_n105, B => 
                           mult_42_I11_n118, CO => mult_42_I11_n65, S => 
                           mult_42_I11_n66);
   mult_42_I11_U43 : FA_X1 port map( A => mult_42_I11_n126, B => 
                           mult_42_I11_n134, CI => mult_42_I11_n142, CO => 
                           mult_42_I11_n63, S => mult_42_I11_n64);
   mult_42_I11_U42 : FA_X1 port map( A => mult_42_I11_n66, B => 
                           mult_42_I11_n151, CI => mult_42_I11_n71, CO => 
                           mult_42_I11_n61, S => mult_42_I11_n62);
   mult_42_I11_U41 : FA_X1 port map( A => mult_42_I11_n64, B => mult_42_I11_n69
                           , CI => mult_42_I11_n62, CO => mult_42_I11_n59, S =>
                           mult_42_I11_n60);
   mult_42_I11_U38 : FA_X1 port map( A => mult_42_I11_n133, B => 
                           mult_42_I11_n117, CI => mult_42_I11_n295, CO => 
                           mult_42_I11_n55, S => mult_42_I11_n56);
   mult_42_I11_U37 : FA_X1 port map( A => mult_42_I11_n58, B => mult_42_I11_n65
                           , CI => mult_42_I11_n63, CO => mult_42_I11_n53, S =>
                           mult_42_I11_n54);
   mult_42_I11_U36 : FA_X1 port map( A => mult_42_I11_n61, B => mult_42_I11_n56
                           , CI => mult_42_I11_n54, CO => mult_42_I11_n51, S =>
                           mult_42_I11_n52);
   mult_42_I11_U34 : FA_X1 port map( A => mult_42_I11_n124, B => 
                           mult_42_I11_n116, CI => mult_42_I11_n132, CO => 
                           mult_42_I11_n47, S => mult_42_I11_n48);
   mult_42_I11_U33 : FA_X1 port map( A => mult_42_I11_n57, B => mult_42_I11_n50
                           , CI => mult_42_I11_n55, CO => mult_42_I11_n45, S =>
                           mult_42_I11_n46);
   mult_42_I11_U32 : FA_X1 port map( A => mult_42_I11_n53, B => mult_42_I11_n48
                           , CI => mult_42_I11_n46, CO => mult_42_I11_n43, S =>
                           mult_42_I11_n44);
   mult_42_I11_U31 : FA_X1 port map( A => mult_42_I11_n123, B => 
                           mult_42_I11_n115, CI => mult_42_I11_n140, CO => 
                           mult_42_I11_n41, S => mult_42_I11_n42);
   mult_42_I11_U30 : FA_X1 port map( A => mult_42_I11_n297, B => 
                           mult_42_I11_n131, CI => mult_42_I11_n47, CO => 
                           mult_42_I11_n39, S => mult_42_I11_n40);
   mult_42_I11_U29 : FA_X1 port map( A => mult_42_I11_n45, B => mult_42_I11_n42
                           , CI => mult_42_I11_n40, CO => mult_42_I11_n37, S =>
                           mult_42_I11_n38);
   mult_42_I11_U27 : FA_X1 port map( A => mult_42_I11_n114, B => 
                           mult_42_I11_n122, CI => mult_42_I11_n299, CO => 
                           mult_42_I11_n33, S => mult_42_I11_n34);
   mult_42_I11_U26 : FA_X1 port map( A => mult_42_I11_n34, B => mult_42_I11_n41
                           , CI => mult_42_I11_n39, CO => mult_42_I11_n31, S =>
                           mult_42_I11_n32);
   mult_42_I11_U25 : FA_X1 port map( A => mult_42_I11_n121, B => 
                           mult_42_I11_n35, CI => mult_42_I11_n298, CO => 
                           mult_42_I11_n29, S => mult_42_I11_n30);
   mult_42_I11_U24 : FA_X1 port map( A => mult_42_I11_n33, B => 
                           mult_42_I11_n113, CI => mult_42_I11_n30, CO => 
                           mult_42_I11_n27, S => mult_42_I11_n28);
   mult_42_I11_U22 : FA_X1 port map( A => mult_42_I11_n301, B => 
                           mult_42_I11_n112, CI => mult_42_I11_n29, CO => 
                           mult_42_I11_n23, S => mult_42_I11_n24);
   mult_42_I11_U21 : FA_X1 port map( A => mult_42_I11_n111, B => 
                           mult_42_I11_n25, CI => mult_42_I11_n300, CO => 
                           mult_42_I11_n21, S => mult_42_I11_n22);
   mult_42_I11_U10 : FA_X1 port map( A => mult_42_I11_n52, B => mult_42_I11_n59
                           , CI => mult_42_I11_n10, CO => mult_42_I11_n9, S => 
                           N193_port);
   mult_42_I11_U9 : FA_X1 port map( A => mult_42_I11_n44, B => mult_42_I11_n51,
                           CI => mult_42_I11_n9, CO => mult_42_I11_n8, S => 
                           N194_port);
   mult_42_I11_U8 : FA_X1 port map( A => mult_42_I11_n38, B => mult_42_I11_n43,
                           CI => mult_42_I11_n8, CO => mult_42_I11_n7, S => 
                           N195_port);
   mult_42_I11_U7 : FA_X1 port map( A => mult_42_I11_n32, B => mult_42_I11_n37,
                           CI => mult_42_I11_n7, CO => mult_42_I11_n6, S => 
                           N196_port);
   mult_42_I11_U6 : FA_X1 port map( A => mult_42_I11_n28, B => mult_42_I11_n31,
                           CI => mult_42_I11_n6, CO => mult_42_I11_n5, S => 
                           N197_port);
   mult_42_I11_U5 : FA_X1 port map( A => mult_42_I11_n24, B => mult_42_I11_n27,
                           CI => mult_42_I11_n5, CO => mult_42_I11_n4, S => 
                           N198_port);
   mult_42_I11_U4 : FA_X1 port map( A => mult_42_I11_n23, B => mult_42_I11_n22,
                           CI => mult_42_I11_n4, CO => mult_42_I11_n3, S => 
                           N199_port);
   mult_42_I11_U3 : FA_X1 port map( A => mult_42_I11_n21, B => mult_42_I11_n303
                           , CI => mult_42_I11_n3, CO => mult_42_I11_n2, S => 
                           N200_port);
   mult_42_I11_U2 : FA_X1 port map( A => mult_42_I11_n302, B => mult_42_I11_n19
                           , CI => mult_42_I11_n2, CO => mult_42_I11_n1, S => 
                           N201_port);
   add_6_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N73, B => N153,
                           Z => N23_port);
   add_6_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N73, A2 => 
                           N153, ZN => add_6_root_add_0_root_add_44_I11_n1);
   add_6_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N154, B => N74,
                           CI => add_6_root_add_0_root_add_44_I11_n1, CO => 
                           add_6_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N24);
   add_6_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N155, B => N75,
                           CI => add_6_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_6_root_add_0_root_add_44_I11_carry_3_port,
                           S => N25);
   add_6_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N156_port, B =>
                           N76, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_3_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_4_port, S => 
                           N26);
   add_6_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N157_port, B =>
                           N77, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_4_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_5_port, S => 
                           N27);
   add_6_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N158_port, B =>
                           N78, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_5_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_6_port, S => 
                           N28);
   add_6_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N159_port, B =>
                           N79, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_6_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_7_port, S => 
                           N29);
   add_6_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N160_port, B =>
                           N80, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_7_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_8_port, S => 
                           N30);
   add_6_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N161_port, B =>
                           N81, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_6_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N31);
   add_6_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N162_port, B =>
                           N82, CI => 
                           add_6_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_6_root_add_0_root_add_44_I11_n_1112, S => N32);
   add_8_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N53, B => N93, 
                           Z => N43);
   add_8_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N53, A2 => N93
                           , ZN => add_8_root_add_0_root_add_44_I11_n1);
   add_8_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N94, B => N54, 
                           CI => add_8_root_add_0_root_add_44_I11_n1, CO => 
                           add_8_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N44);
   add_8_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N95, B => N55, 
                           CI => add_8_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_3_port,
                           S => N45);
   add_8_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N96, B => N56, 
                           CI => add_8_root_add_0_root_add_44_I11_carry_3_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_4_port,
                           S => N46);
   add_8_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N97, B => N57, 
                           CI => add_8_root_add_0_root_add_44_I11_carry_4_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_5_port,
                           S => N47);
   add_8_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N98, B => N58, 
                           CI => add_8_root_add_0_root_add_44_I11_carry_5_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_6_port,
                           S => N48);
   add_8_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N99, B => N59, 
                           CI => add_8_root_add_0_root_add_44_I11_carry_6_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_7_port,
                           S => N49);
   add_8_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N100, B => N60,
                           CI => add_8_root_add_0_root_add_44_I11_carry_7_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_8_port,
                           S => N50);
   add_8_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N101, B => N61,
                           CI => add_8_root_add_0_root_add_44_I11_carry_8_port,
                           CO => add_8_root_add_0_root_add_44_I11_carry_9_port,
                           S => N51);
   add_8_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N102, B => N62,
                           CI => add_8_root_add_0_root_add_44_I11_carry_9_port,
                           CO => add_8_root_add_0_root_add_44_I11_n_1115, S => 
                           N52);
   add_9_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N173_port, B =>
                           N133, Z => N63);
   add_9_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N173_port, A2 
                           => N133, ZN => add_9_root_add_0_root_add_44_I11_n1);
   add_9_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N134, B => 
                           N174_port, CI => add_9_root_add_0_root_add_44_I11_n1
                           , CO => 
                           add_9_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N64);
   add_9_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N135, B => 
                           N175_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_2_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_3_port, S => 
                           N65);
   add_9_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N136, B => 
                           N176_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_3_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_4_port, S => 
                           N66);
   add_9_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N137, B => 
                           N177_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_4_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_5_port, S => 
                           N67);
   add_9_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N138, B => 
                           N178_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_5_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_6_port, S => 
                           N68);
   add_9_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N139, B => 
                           N179_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_6_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_7_port, S => 
                           N69);
   add_9_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N140, B => 
                           N180_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_7_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_8_port, S => 
                           N70);
   add_9_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N141, B => 
                           N181_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_9_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N71);
   add_9_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N142, B => 
                           N182_port, CI => 
                           add_9_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_9_root_add_0_root_add_44_I11_n_1118, S => 
                           N72_port);
   add_7_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N113, B => N13,
                           Z => N143);
   add_7_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N113, A2 => 
                           N13, ZN => add_7_root_add_0_root_add_44_I11_n1);
   add_7_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N14, B => N114,
                           CI => add_7_root_add_0_root_add_44_I11_n1, CO => 
                           add_7_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N144);
   add_7_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N15, B => N115,
                           CI => add_7_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_3_port,
                           S => N145);
   add_7_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N16, B => N116,
                           CI => add_7_root_add_0_root_add_44_I11_carry_3_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_4_port,
                           S => N146);
   add_7_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N17, B => N117,
                           CI => add_7_root_add_0_root_add_44_I11_carry_4_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_5_port,
                           S => N147);
   add_7_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N18, B => N118,
                           CI => add_7_root_add_0_root_add_44_I11_carry_5_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_6_port,
                           S => N148);
   add_7_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N19, B => N119,
                           CI => add_7_root_add_0_root_add_44_I11_carry_6_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_7_port,
                           S => N149);
   add_7_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N20, B => N120,
                           CI => add_7_root_add_0_root_add_44_I11_carry_7_port,
                           CO => add_7_root_add_0_root_add_44_I11_carry_8_port,
                           S => N150);
   add_7_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N21_port, B => 
                           N121, CI => 
                           add_7_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_7_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N151);
   add_7_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N22, B => N122,
                           CI => add_7_root_add_0_root_add_44_I11_carry_9_port,
                           CO => add_7_root_add_0_root_add_44_I11_n_1121, S => 
                           N152);
   add_2_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N143, B => 
                           N23_port, Z => N83);
   add_2_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N143, A2 => 
                           N23_port, ZN => add_2_root_add_0_root_add_44_I11_n1)
                           ;
   add_2_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N24, B => N144,
                           CI => add_2_root_add_0_root_add_44_I11_n1, CO => 
                           add_2_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N84);
   add_2_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N25, B => N145,
                           CI => add_2_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_3_port,
                           S => N85);
   add_2_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N26, B => N146,
                           CI => add_2_root_add_0_root_add_44_I11_carry_3_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_4_port,
                           S => N86);
   add_2_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N27, B => N147,
                           CI => add_2_root_add_0_root_add_44_I11_carry_4_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_5_port,
                           S => N87);
   add_2_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N28, B => N148,
                           CI => add_2_root_add_0_root_add_44_I11_carry_5_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_6_port,
                           S => N88);
   add_2_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N29, B => N149,
                           CI => add_2_root_add_0_root_add_44_I11_carry_6_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_7_port,
                           S => N89);
   add_2_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N30, B => N150,
                           CI => add_2_root_add_0_root_add_44_I11_carry_7_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_8_port,
                           S => N90);
   add_2_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N31, B => N151,
                           CI => add_2_root_add_0_root_add_44_I11_carry_8_port,
                           CO => add_2_root_add_0_root_add_44_I11_carry_9_port,
                           S => N91);
   add_2_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N32, B => N152,
                           CI => add_2_root_add_0_root_add_44_I11_carry_9_port,
                           CO => add_2_root_add_0_root_add_44_I11_n_1124, S => 
                           N92);
   add_3_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N63, B => N43, 
                           Z => N103);
   add_3_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N63, A2 => N43
                           , ZN => add_3_root_add_0_root_add_44_I11_n1);
   add_3_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N44, B => N64, 
                           CI => add_3_root_add_0_root_add_44_I11_n1, CO => 
                           add_3_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N104);
   add_3_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N45, B => N65, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_3_port,
                           S => N105);
   add_3_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N46, B => N66, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_3_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_4_port,
                           S => N106);
   add_3_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N47, B => N67, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_4_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_5_port,
                           S => N107);
   add_3_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N48, B => N68, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_5_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_6_port,
                           S => N108);
   add_3_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N49, B => N69, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_6_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_7_port,
                           S => N109);
   add_3_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N50, B => N70, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_7_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_8_port,
                           S => N110);
   add_3_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N51, B => N71, 
                           CI => add_3_root_add_0_root_add_44_I11_carry_8_port,
                           CO => add_3_root_add_0_root_add_44_I11_carry_9_port,
                           S => N111);
   add_3_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N52, B => 
                           N72_port, CI => 
                           add_3_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_3_root_add_0_root_add_44_I11_n_1127, S => N112);
   add_5_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N193_port, B =>
                           N3, Z => N123);
   add_5_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N193_port, A2 
                           => N3, ZN => add_5_root_add_0_root_add_44_I11_n1);
   add_5_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N4, B => 
                           N194_port, CI => add_5_root_add_0_root_add_44_I11_n1
                           , CO => 
                           add_5_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N124);
   add_5_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N5, B => 
                           N195_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_2_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_3_port, S => 
                           N125);
   add_5_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N6, B => 
                           N196_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_3_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_4_port, S => 
                           N126);
   add_5_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N7, B => 
                           N197_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_4_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_5_port, S => 
                           N127);
   add_5_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N8, B => 
                           N198_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_5_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_6_port, S => 
                           N128);
   add_5_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N9, B => 
                           N199_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_6_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_7_port, S => 
                           N129);
   add_5_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N10, B => 
                           N200_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_7_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_8_port, S => 
                           N130);
   add_5_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N11, B => 
                           N201_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_5_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N131);
   add_5_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N12, B => 
                           N202_port, CI => 
                           add_5_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_5_root_add_0_root_add_44_I11_n_1130, S => N132);
   add_4_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N123, B => N33,
                           Z => N183_port);
   add_4_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N123, A2 => 
                           N33, ZN => add_4_root_add_0_root_add_44_I11_n1);
   add_4_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N34, B => N124,
                           CI => add_4_root_add_0_root_add_44_I11_n1, CO => 
                           add_4_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N184_port);
   add_4_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N35, B => N125,
                           CI => add_4_root_add_0_root_add_44_I11_carry_2_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_3_port,
                           S => N185_port);
   add_4_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N36, B => N126,
                           CI => add_4_root_add_0_root_add_44_I11_carry_3_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_4_port,
                           S => N186_port);
   add_4_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N37, B => N127,
                           CI => add_4_root_add_0_root_add_44_I11_carry_4_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_5_port,
                           S => N187_port);
   add_4_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N38, B => N128,
                           CI => add_4_root_add_0_root_add_44_I11_carry_5_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_6_port,
                           S => N188_port);
   add_4_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N39, B => N129,
                           CI => add_4_root_add_0_root_add_44_I11_carry_6_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_7_port,
                           S => N189_port);
   add_4_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N40, B => N130,
                           CI => add_4_root_add_0_root_add_44_I11_carry_7_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_8_port,
                           S => N190_port);
   add_4_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N41, B => N131,
                           CI => add_4_root_add_0_root_add_44_I11_carry_8_port,
                           CO => add_4_root_add_0_root_add_44_I11_carry_9_port,
                           S => N191_port);
   add_4_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N42, B => N132,
                           CI => add_4_root_add_0_root_add_44_I11_carry_9_port,
                           CO => add_4_root_add_0_root_add_44_I11_n_1133, S => 
                           N192_port);
   add_1_root_add_0_root_add_44_I11_U2 : XOR2_X1 port map( A => N83, B => 
                           N183_port, Z => N163_port);
   add_1_root_add_0_root_add_44_I11_U1 : AND2_X1 port map( A1 => N83, A2 => 
                           N183_port, ZN => add_1_root_add_0_root_add_44_I11_n1
                           );
   add_1_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N184_port, B =>
                           N84, CI => add_1_root_add_0_root_add_44_I11_n1, CO 
                           => add_1_root_add_0_root_add_44_I11_carry_2_port, S 
                           => N164_port);
   add_1_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N185_port, B =>
                           N85, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_2_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_3_port, S => 
                           N165_port);
   add_1_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N186_port, B =>
                           N86, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_3_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_4_port, S => 
                           N166_port);
   add_1_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N187_port, B =>
                           N87, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_4_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_5_port, S => 
                           N167_port);
   add_1_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N188_port, B =>
                           N88, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_5_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_6_port, S => 
                           N168_port);
   add_1_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N189_port, B =>
                           N89, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_6_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_7_port, S => 
                           N169_port);
   add_1_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N190_port, B =>
                           N90, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_7_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_8_port, S => 
                           N170_port);
   add_1_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N191_port, B =>
                           N91, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_1_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N171_port);
   add_1_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N192_port, B =>
                           N92, CI => 
                           add_1_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_1_root_add_0_root_add_44_I11_n_1136, S => 
                           N172_port);
   add_0_root_add_0_root_add_44_I11_U2 : AND2_X1 port map( A1 => N163_port, A2 
                           => N103, ZN => add_0_root_add_0_root_add_44_I11_n2);
   add_0_root_add_0_root_add_44_I11_U1 : XOR2_X1 port map( A => N163_port, B =>
                           N103, Z => N203);
   add_0_root_add_0_root_add_44_I11_U1_1 : FA_X1 port map( A => N104, B => 
                           N164_port, CI => add_0_root_add_0_root_add_44_I11_n2
                           , CO => 
                           add_0_root_add_0_root_add_44_I11_carry_2_port, S => 
                           N204);
   add_0_root_add_0_root_add_44_I11_U1_2 : FA_X1 port map( A => N105, B => 
                           N165_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_2_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_3_port, S => 
                           N205);
   add_0_root_add_0_root_add_44_I11_U1_3 : FA_X1 port map( A => N106, B => 
                           N166_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_3_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_4_port, S => 
                           N206);
   add_0_root_add_0_root_add_44_I11_U1_4 : FA_X1 port map( A => N107, B => 
                           N167_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_4_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_5_port, S => 
                           N207);
   add_0_root_add_0_root_add_44_I11_U1_5 : FA_X1 port map( A => N108, B => 
                           N168_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_5_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_6_port, S => 
                           N208);
   add_0_root_add_0_root_add_44_I11_U1_6 : FA_X1 port map( A => N109, B => 
                           N169_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_6_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_7_port, S => 
                           N209);
   add_0_root_add_0_root_add_44_I11_U1_7 : FA_X1 port map( A => N110, B => 
                           N170_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_7_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_8_port, S => 
                           N210);
   add_0_root_add_0_root_add_44_I11_U1_8 : FA_X1 port map( A => N111, B => 
                           N171_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_8_port, CO =>
                           add_0_root_add_0_root_add_44_I11_carry_9_port, S => 
                           N211);
   add_0_root_add_0_root_add_44_I11_U1_9 : FA_X1 port map( A => N112, B => 
                           N172_port, CI => 
                           add_0_root_add_0_root_add_44_I11_carry_9_port, CO =>
                           add_0_root_add_0_root_add_44_I11_n_1139, S => N212);

end SYN_beh;
